.SUBCKT CIM rst_n clk in_valid weight_valid out_valid Out_OFM[12] Out_OFM[11] Out_OFM[10] Out_OFM[9] Out_OFM[8] Out_OFM[7] Out_OFM[6] Out_OFM[5] Out_OFM[4] Out_OFM[3] Out_OFM[2] Out_OFM[1] Out_OFM[0]
Xclk21_reg n1269 clk n1905 n1254 clk21 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM1_reg_12_ n680 n1269 Out_OFM1[12] DFFHQNx1_ASAP7_75t_R
XOut_OFM1_reg_11_ n679 n1269 Out_OFM1[11] DFFHQNx1_ASAP7_75t_R
XOut_OFM1_reg_10_ n678 n1269 Out_OFM1[10] DFFHQNx1_ASAP7_75t_R
XOut_OFM1_reg_9_ n677 n1269 Out_OFM1[9] DFFHQNx1_ASAP7_75t_R
XOut_OFM1_reg_8_ n676 n1269 Out_OFM1[8] DFFHQNx1_ASAP7_75t_R
XOut_OFM1_reg_7_ n675 n1269 Out_OFM1[7] DFFHQNx1_ASAP7_75t_R
XOut_OFM1_reg_6_ n674 n1269 Out_OFM1[6] DFFHQNx1_ASAP7_75t_R
XOut_OFM1_reg_5_ n673 n1269 Out_OFM1[5] DFFHQNx1_ASAP7_75t_R
XOut_OFM1_reg_4_ n672 n1269 Out_OFM1[4] DFFHQNx1_ASAP7_75t_R
XOut_OFM1_reg_3_ n671 n1269 Out_OFM1[3] DFFHQNx1_ASAP7_75t_R
XOut_OFM1_reg_2_ n670 n1269 Out_OFM1[2] DFFHQNx1_ASAP7_75t_R
XOut_OFM1_reg_1_ n669 n1269 Out_OFM1[1] DFFHQNx1_ASAP7_75t_R
XOut_OFM1_reg_0_ n668 n1269 Out_OFM1[0] DFFHQNx1_ASAP7_75t_R
XOut_OFM2_reg_12_ n680 clk22 Out_OFM2[12] DFFHQNx1_ASAP7_75t_R
XOut_OFM2_reg_11_ n679 clk22 Out_OFM2[11] DFFHQNx1_ASAP7_75t_R
XOut_OFM2_reg_10_ n678 clk22 Out_OFM2[10] DFFHQNx1_ASAP7_75t_R
XOut_OFM2_reg_9_ n677 clk22 Out_OFM2[9] DFFHQNx1_ASAP7_75t_R
XOut_OFM2_reg_8_ n676 clk22 Out_OFM2[8] DFFHQNx1_ASAP7_75t_R
XOut_OFM2_reg_7_ n675 clk22 Out_OFM2[7] DFFHQNx1_ASAP7_75t_R
XOut_OFM2_reg_6_ n674 clk22 Out_OFM2[6] DFFHQNx1_ASAP7_75t_R
XOut_OFM2_reg_5_ n673 clk22 Out_OFM2[5] DFFHQNx1_ASAP7_75t_R
XOut_OFM2_reg_4_ n672 clk22 Out_OFM2[4] DFFHQNx1_ASAP7_75t_R
XOut_OFM2_reg_3_ n671 clk22 Out_OFM2[3] DFFHQNx1_ASAP7_75t_R
XOut_OFM2_reg_2_ n670 clk22 Out_OFM2[2] DFFHQNx1_ASAP7_75t_R
XOut_OFM2_reg_1_ n669 clk22 Out_OFM2[1] DFFHQNx1_ASAP7_75t_R
XOut_OFM2_reg_0_ n668 clk22 Out_OFM2[0] DFFHQNx1_ASAP7_75t_R
XU17 n125 n126 n681 OR2x2_ASAP7_75t_R
XU20 n128 n129 n683 OR2x2_ASAP7_75t_R
XU23 n130 n131 n685 OR2x2_ASAP7_75t_R
XU26 n132 n133 n687 OR2x2_ASAP7_75t_R
XU29 n134 n135 n689 OR2x2_ASAP7_75t_R
XU32 n136 n137 n691 OR2x2_ASAP7_75t_R
XU35 n138 n139 n693 OR2x2_ASAP7_75t_R
XU38 n140 n141 n695 OR2x2_ASAP7_75t_R
XU41 n142 n143 n697 OR2x2_ASAP7_75t_R
XU44 n144 n145 n699 OR2x2_ASAP7_75t_R
XU47 n146 n147 n701 OR2x2_ASAP7_75t_R
XU50 n148 n149 n703 OR2x2_ASAP7_75t_R
XU53 n150 n151 n705 OR2x2_ASAP7_75t_R
XU56 n152 n153 n707 OR2x2_ASAP7_75t_R
XU59 n154 n155 n709 OR2x2_ASAP7_75t_R
XU62 n156 n157 n711 OR2x2_ASAP7_75t_R
XU65 n158 n159 n713 OR2x2_ASAP7_75t_R
XU68 n160 n161 n715 OR2x2_ASAP7_75t_R
XU71 n162 n163 n717 OR2x2_ASAP7_75t_R
XU74 n164 n165 n719 OR2x2_ASAP7_75t_R
XU77 n166 n167 n721 OR2x2_ASAP7_75t_R
XU80 n168 n169 n723 OR2x2_ASAP7_75t_R
XU83 n170 n171 n725 OR2x2_ASAP7_75t_R
XU86 n172 n173 n727 OR2x2_ASAP7_75t_R
XU89 n174 n175 n729 OR2x2_ASAP7_75t_R
XU92 n176 n177 n731 OR2x2_ASAP7_75t_R
XU95 n178 n179 n733 OR2x2_ASAP7_75t_R
XU98 n180 n181 n735 OR2x2_ASAP7_75t_R
XU101 n182 n183 n737 OR2x2_ASAP7_75t_R
XU104 n184 n185 n739 OR2x2_ASAP7_75t_R
XU107 n186 n187 n741 OR2x2_ASAP7_75t_R
XU110 n188 n189 n743 OR2x2_ASAP7_75t_R
XU113 n190 n191 n745 OR2x2_ASAP7_75t_R
XU116 n192 n193 n747 OR2x2_ASAP7_75t_R
XU119 n194 n195 n749 OR2x2_ASAP7_75t_R
XU122 n196 n197 n751 OR2x2_ASAP7_75t_R
XU125 n198 n199 n753 OR2x2_ASAP7_75t_R
XU128 n200 n201 n755 OR2x2_ASAP7_75t_R
XU131 n202 n203 n757 OR2x2_ASAP7_75t_R
XU134 n204 n205 n759 OR2x2_ASAP7_75t_R
XU137 n206 n207 n761 OR2x2_ASAP7_75t_R
XU140 n208 n209 n763 OR2x2_ASAP7_75t_R
XU143 n210 n211 n765 OR2x2_ASAP7_75t_R
XU146 n212 n213 n767 OR2x2_ASAP7_75t_R
XU149 n214 n215 n769 OR2x2_ASAP7_75t_R
XU152 n216 n217 n771 OR2x2_ASAP7_75t_R
XU155 n218 n219 n773 OR2x2_ASAP7_75t_R
XU158 n220 n221 n775 OR2x2_ASAP7_75t_R
XU161 n222 n223 n777 OR2x2_ASAP7_75t_R
XU164 n224 n225 n779 OR2x2_ASAP7_75t_R
XU167 n226 n227 n781 OR2x2_ASAP7_75t_R
XU170 n228 n229 n783 OR2x2_ASAP7_75t_R
XU173 n230 n231 n785 OR2x2_ASAP7_75t_R
XU176 n232 n233 n787 OR2x2_ASAP7_75t_R
XU179 n234 n235 n789 OR2x2_ASAP7_75t_R
XU182 n236 n237 n791 OR2x2_ASAP7_75t_R
XU185 n238 n239 n793 OR2x2_ASAP7_75t_R
XU188 n240 n241 n795 OR2x2_ASAP7_75t_R
XU191 n242 n243 n797 OR2x2_ASAP7_75t_R
XU194 n244 n245 n799 OR2x2_ASAP7_75t_R
XU197 n246 n247 n801 OR2x2_ASAP7_75t_R
XU200 n248 n249 n803 OR2x2_ASAP7_75t_R
XU203 n250 n251 n805 OR2x2_ASAP7_75t_R
XU206 n252 n253 n807 OR2x2_ASAP7_75t_R
XU209 n254 n255 n809 OR2x2_ASAP7_75t_R
XU212 n256 n257 n811 OR2x2_ASAP7_75t_R
XU215 n258 n259 n813 OR2x2_ASAP7_75t_R
XU218 n260 n261 n815 OR2x2_ASAP7_75t_R
XU221 n262 n263 n817 OR2x2_ASAP7_75t_R
XU224 n264 n265 n819 OR2x2_ASAP7_75t_R
XU227 n266 n267 n821 OR2x2_ASAP7_75t_R
XU230 n268 n269 n823 OR2x2_ASAP7_75t_R
XU233 n270 n271 n825 OR2x2_ASAP7_75t_R
XU236 n272 n273 n827 OR2x2_ASAP7_75t_R
XU239 n274 n275 n829 OR2x2_ASAP7_75t_R
XU242 n276 n277 n831 OR2x2_ASAP7_75t_R
XU245 n278 n279 n833 OR2x2_ASAP7_75t_R
XU248 n280 n281 n835 OR2x2_ASAP7_75t_R
XU251 n282 n283 n837 OR2x2_ASAP7_75t_R
XU254 n284 n285 n839 OR2x2_ASAP7_75t_R
XU257 n286 n287 n841 OR2x2_ASAP7_75t_R
XU260 n288 n289 n843 OR2x2_ASAP7_75t_R
XU263 n290 n291 n845 OR2x2_ASAP7_75t_R
XU266 n292 n293 n847 OR2x2_ASAP7_75t_R
XU269 n294 n295 n849 OR2x2_ASAP7_75t_R
XU272 n296 n297 n851 OR2x2_ASAP7_75t_R
XU275 n298 n299 n853 OR2x2_ASAP7_75t_R
XU278 n300 n301 n855 OR2x2_ASAP7_75t_R
XU281 n302 n303 n857 OR2x2_ASAP7_75t_R
XU284 n304 n305 n859 OR2x2_ASAP7_75t_R
XU287 n306 n307 n861 OR2x2_ASAP7_75t_R
XU290 n308 n309 n863 OR2x2_ASAP7_75t_R
XU293 n310 n311 n865 OR2x2_ASAP7_75t_R
XU296 n312 n313 n867 OR2x2_ASAP7_75t_R
XU299 n314 n315 n869 OR2x2_ASAP7_75t_R
XU302 n316 n317 n871 OR2x2_ASAP7_75t_R
XU305 n318 n319 n873 OR2x2_ASAP7_75t_R
XU308 n320 n321 n875 OR2x2_ASAP7_75t_R
XU311 n322 n323 n877 OR2x2_ASAP7_75t_R
XU314 n324 n325 n879 OR2x2_ASAP7_75t_R
XU317 n326 n327 n881 OR2x2_ASAP7_75t_R
XU320 n328 n329 n883 OR2x2_ASAP7_75t_R
XU323 n330 n331 n885 OR2x2_ASAP7_75t_R
XU326 n332 n333 n887 OR2x2_ASAP7_75t_R
XU329 n334 n335 n889 OR2x2_ASAP7_75t_R
XU332 n336 n337 n891 OR2x2_ASAP7_75t_R
XU335 n338 n339 n893 OR2x2_ASAP7_75t_R
XU338 n340 n341 n895 OR2x2_ASAP7_75t_R
XU341 n342 n343 n897 OR2x2_ASAP7_75t_R
XU344 n344 n345 n899 OR2x2_ASAP7_75t_R
XU347 n346 n347 n901 OR2x2_ASAP7_75t_R
XU350 n348 n349 n903 OR2x2_ASAP7_75t_R
XU353 n350 n351 n905 OR2x2_ASAP7_75t_R
XU356 n352 n353 n907 OR2x2_ASAP7_75t_R
XU359 n354 n355 n909 OR2x2_ASAP7_75t_R
XU362 n356 n357 n911 OR2x2_ASAP7_75t_R
XU365 n358 n359 n913 OR2x2_ASAP7_75t_R
XU368 n360 n361 n915 OR2x2_ASAP7_75t_R
XU371 n362 n363 n917 OR2x2_ASAP7_75t_R
XU374 n364 n365 n919 OR2x2_ASAP7_75t_R
XU377 n366 n367 n921 OR2x2_ASAP7_75t_R
XU380 n368 n369 n923 OR2x2_ASAP7_75t_R
XU383 n370 n371 n925 OR2x2_ASAP7_75t_R
XU386 n372 n373 n927 OR2x2_ASAP7_75t_R
XU389 n374 n375 n929 OR2x2_ASAP7_75t_R
XU392 n376 n377 n931 OR2x2_ASAP7_75t_R
XU395 n378 n379 n933 OR2x2_ASAP7_75t_R
XU398 n380 n381 n935 OR2x2_ASAP7_75t_R
XU402 n382 n383 n937 OR2x2_ASAP7_75t_R
XU405 n384 n385 n939 OR2x2_ASAP7_75t_R
XU408 n386 n387 n941 OR2x2_ASAP7_75t_R
XU411 n388 n389 n943 OR2x2_ASAP7_75t_R
XU414 n390 n391 n945 OR2x2_ASAP7_75t_R
XU417 n392 n393 n947 OR2x2_ASAP7_75t_R
XU420 n394 n395 n949 OR2x2_ASAP7_75t_R
XU423 n396 n397 n951 OR2x2_ASAP7_75t_R
XU426 n398 n399 n953 OR2x2_ASAP7_75t_R
XU429 n400 n401 n955 OR2x2_ASAP7_75t_R
XU432 n402 n403 n957 OR2x2_ASAP7_75t_R
XU435 n404 n405 n959 OR2x2_ASAP7_75t_R
XU438 n406 n407 n961 OR2x2_ASAP7_75t_R
XU441 n408 n409 n963 OR2x2_ASAP7_75t_R
XU444 n410 n411 n965 OR2x2_ASAP7_75t_R
XU447 n412 n413 n967 OR2x2_ASAP7_75t_R
XU450 n414 n415 n969 OR2x2_ASAP7_75t_R
XU453 n416 n417 n971 OR2x2_ASAP7_75t_R
XU456 n418 n419 n973 OR2x2_ASAP7_75t_R
XU459 n420 n421 n975 OR2x2_ASAP7_75t_R
XU462 n422 n423 n977 OR2x2_ASAP7_75t_R
XU465 n424 n425 n979 OR2x2_ASAP7_75t_R
XU468 n426 n427 n981 OR2x2_ASAP7_75t_R
XU471 n428 n429 n983 OR2x2_ASAP7_75t_R
XU474 n430 n431 n985 OR2x2_ASAP7_75t_R
XU477 n432 n433 n987 OR2x2_ASAP7_75t_R
XU480 n434 n435 n989 OR2x2_ASAP7_75t_R
XU483 n436 n437 n991 OR2x2_ASAP7_75t_R
XU486 n438 n439 n993 OR2x2_ASAP7_75t_R
XU489 n440 n441 n995 OR2x2_ASAP7_75t_R
XU492 n442 n443 n997 OR2x2_ASAP7_75t_R
XU495 n444 n445 n999 OR2x2_ASAP7_75t_R
XU498 n446 n447 n1001 OR2x2_ASAP7_75t_R
XU501 n448 n449 n1003 OR2x2_ASAP7_75t_R
XU504 n450 n451 n1005 OR2x2_ASAP7_75t_R
XU507 n452 n453 n1007 OR2x2_ASAP7_75t_R
XU510 n454 n455 n1009 OR2x2_ASAP7_75t_R
XU513 n456 n457 n1011 OR2x2_ASAP7_75t_R
XU516 n458 n459 n1013 OR2x2_ASAP7_75t_R
XU519 n460 n461 n1015 OR2x2_ASAP7_75t_R
XU522 n462 n463 n1017 OR2x2_ASAP7_75t_R
XU525 n464 n465 n1019 OR2x2_ASAP7_75t_R
XU528 n466 n467 n1021 OR2x2_ASAP7_75t_R
XU531 n468 n469 n1023 OR2x2_ASAP7_75t_R
XU534 n470 n471 n1025 OR2x2_ASAP7_75t_R
XU537 n472 n473 n1027 OR2x2_ASAP7_75t_R
XU540 n474 n475 n1029 OR2x2_ASAP7_75t_R
XU543 n476 n477 n1031 OR2x2_ASAP7_75t_R
XU546 n478 n479 n1033 OR2x2_ASAP7_75t_R
XU549 n480 n481 n1035 OR2x2_ASAP7_75t_R
XU552 n482 n483 n1037 OR2x2_ASAP7_75t_R
XU555 n484 n485 n1039 OR2x2_ASAP7_75t_R
XU558 n486 n487 n1041 OR2x2_ASAP7_75t_R
XU561 n488 n489 n1043 OR2x2_ASAP7_75t_R
XU564 n490 n491 n1045 OR2x2_ASAP7_75t_R
XU567 n492 n493 n1047 OR2x2_ASAP7_75t_R
XU570 n494 n495 n1049 OR2x2_ASAP7_75t_R
XU573 n496 n497 n1051 OR2x2_ASAP7_75t_R
XU576 n498 n499 n1053 OR2x2_ASAP7_75t_R
XU579 n500 n501 n1055 OR2x2_ASAP7_75t_R
XU582 n502 n503 n1057 OR2x2_ASAP7_75t_R
XU585 n504 n505 n1059 OR2x2_ASAP7_75t_R
XU588 n506 n507 n1061 OR2x2_ASAP7_75t_R
XU591 n508 n509 n1063 OR2x2_ASAP7_75t_R
XU594 n510 n511 n1065 OR2x2_ASAP7_75t_R
XU597 n512 n513 n1067 OR2x2_ASAP7_75t_R
XU600 n514 n515 n1069 OR2x2_ASAP7_75t_R
XU603 n516 n517 n1071 OR2x2_ASAP7_75t_R
XU606 n518 n519 n1073 OR2x2_ASAP7_75t_R
XU609 n520 n521 n1075 OR2x2_ASAP7_75t_R
XU612 n522 n523 n1077 OR2x2_ASAP7_75t_R
XU615 n524 n525 n1079 OR2x2_ASAP7_75t_R
XU618 n526 n527 n1081 OR2x2_ASAP7_75t_R
XU621 n528 n529 n1083 OR2x2_ASAP7_75t_R
XU624 n530 n531 n1085 OR2x2_ASAP7_75t_R
XU627 n532 n533 n1087 OR2x2_ASAP7_75t_R
XU630 n534 n535 n1089 OR2x2_ASAP7_75t_R
XU633 n536 n537 n1091 OR2x2_ASAP7_75t_R
XU636 n538 n539 n1093 OR2x2_ASAP7_75t_R
XU639 n540 n541 n1095 OR2x2_ASAP7_75t_R
XU642 n542 n543 n1097 OR2x2_ASAP7_75t_R
XU645 n544 n545 n1099 OR2x2_ASAP7_75t_R
XU648 n546 n547 n1101 OR2x2_ASAP7_75t_R
XU651 n548 n549 n1103 OR2x2_ASAP7_75t_R
XU654 n550 n551 n1105 OR2x2_ASAP7_75t_R
XU657 n552 n553 n1107 OR2x2_ASAP7_75t_R
XU660 n554 n555 n1109 OR2x2_ASAP7_75t_R
XU663 n556 n557 n1111 OR2x2_ASAP7_75t_R
XU666 n558 n559 n1113 OR2x2_ASAP7_75t_R
XU669 n560 n561 n1115 OR2x2_ASAP7_75t_R
XU672 n562 n563 n1117 OR2x2_ASAP7_75t_R
XU675 n564 n565 n1119 OR2x2_ASAP7_75t_R
XU678 n566 n567 n1121 OR2x2_ASAP7_75t_R
XU681 n568 n569 n1123 OR2x2_ASAP7_75t_R
XU684 n570 n571 n1125 OR2x2_ASAP7_75t_R
XU687 n572 n573 n1127 OR2x2_ASAP7_75t_R
XU690 n574 n575 n1129 OR2x2_ASAP7_75t_R
XU693 n576 n577 n1131 OR2x2_ASAP7_75t_R
XU696 n578 n579 n1133 OR2x2_ASAP7_75t_R
XU699 n580 n581 n1135 OR2x2_ASAP7_75t_R
XU702 n582 n583 n1137 OR2x2_ASAP7_75t_R
XU705 n584 n585 n1139 OR2x2_ASAP7_75t_R
XU708 n586 n587 n1141 OR2x2_ASAP7_75t_R
XU711 n588 n589 n1143 OR2x2_ASAP7_75t_R
XU714 n590 n591 n1145 OR2x2_ASAP7_75t_R
XU717 n592 n593 n1147 OR2x2_ASAP7_75t_R
XU720 n594 n595 n1149 OR2x2_ASAP7_75t_R
XU723 n596 n597 n1151 OR2x2_ASAP7_75t_R
XU726 n598 n599 n1153 OR2x2_ASAP7_75t_R
XU729 n600 n601 n1155 OR2x2_ASAP7_75t_R
XU732 n602 n603 n1157 OR2x2_ASAP7_75t_R
XU735 n604 n605 n1159 OR2x2_ASAP7_75t_R
XU738 n606 n607 n1161 OR2x2_ASAP7_75t_R
XU741 n608 n609 n1163 OR2x2_ASAP7_75t_R
XU744 n610 n611 n1165 OR2x2_ASAP7_75t_R
XU747 n612 n613 n1167 OR2x2_ASAP7_75t_R
XU750 n614 n615 n1169 OR2x2_ASAP7_75t_R
XU753 n616 n617 n1171 OR2x2_ASAP7_75t_R
XU756 n618 n619 n1173 OR2x2_ASAP7_75t_R
XU759 n620 n621 n1175 OR2x2_ASAP7_75t_R
XU762 n622 n623 n1177 OR2x2_ASAP7_75t_R
XU765 n624 n625 n1179 OR2x2_ASAP7_75t_R
XU768 n626 n627 n1181 OR2x2_ASAP7_75t_R
XU771 n628 n629 n1183 OR2x2_ASAP7_75t_R
XU774 n630 n631 n1185 OR2x2_ASAP7_75t_R
XU777 n632 n633 n1187 OR2x2_ASAP7_75t_R
XU780 n634 n635 n1189 OR2x2_ASAP7_75t_R
XU783 n636 n637 n1191 OR2x2_ASAP7_75t_R
Xr801 IFM[127] IFM[126] IFM[125] IFM[124] Weight[127] Weight[126] Weight[125] Weight[124] N17 N16 N15 N14 N13 N12 N11 N10 CIM_DW_mult_uns_31
Xr802 IFM[123] IFM[122] IFM[121] IFM[120] Weight[123] Weight[122] Weight[121] Weight[120] N25 N24 N23 N22 N21 N20 N19 N18 CIM_DW_mult_uns_30
Xr804 IFM[119] IFM[118] IFM[117] IFM[116] Weight[119] Weight[118] Weight[117] Weight[116] N704 N703 N702 N701 N700 N699 N698 N697 CIM_DW_mult_uns_29
Xr806 IFM[115] IFM[114] IFM[113] IFM[112] Weight[115] Weight[114] Weight[113] Weight[112] N722 N721 N720 N719 N718 N717 N716 N715 CIM_DW_mult_uns_28
Xr808 IFM[111] IFM[110] IFM[109] IFM[108] Weight[111] Weight[110] Weight[109] Weight[108] N741 N740 N739 N738 N737 N736 N735 N734 CIM_DW_mult_uns_27
Xr810 IFM[107] IFM[106] IFM[105] IFM[104] Weight[107] Weight[106] Weight[105] Weight[104] N761 N760 N759 N758 N757 N756 N755 N754 CIM_DW_mult_uns_26
Xr812 IFM[103] IFM[102] IFM[101] IFM[100] Weight[103] Weight[102] Weight[101] Weight[100] N782 N781 N780 N779 N778 N777 N776 N775 CIM_DW_mult_uns_25
Xr814 IFM[99] IFM[98] IFM[97] IFM[96] Weight[99] Weight[98] Weight[97] Weight[96] N803 N802 N801 N800 N799 N798 N797 N796 CIM_DW_mult_uns_24
Xr816 IFM[95] IFM[94] IFM[93] IFM[92] Weight[95] Weight[94] Weight[93] Weight[92] N824 N823 N822 N821 N820 N819 N818 N817 CIM_DW_mult_uns_23
Xr818 IFM[91] IFM[90] IFM[89] IFM[88] Weight[91] Weight[90] Weight[89] Weight[88] N845 N844 N843 N842 N841 N840 N839 N838 CIM_DW_mult_uns_22
Xr820 IFM[87] IFM[86] IFM[85] IFM[84] Weight[87] Weight[86] Weight[85] Weight[84] N866 N865 N864 N863 N862 N861 N860 N859 CIM_DW_mult_uns_21
Xr822 IFM[83] IFM[82] IFM[81] IFM[80] Weight[83] Weight[82] Weight[81] Weight[80] N887 N886 N885 N884 N883 N882 N881 N880 CIM_DW_mult_uns_20
Xr824 IFM[79] IFM[78] IFM[77] IFM[76] Weight[79] Weight[78] Weight[77] Weight[76] N908 N907 N906 N905 N904 N903 N902 N901 CIM_DW_mult_uns_19
Xr826 IFM[75] IFM[74] IFM[73] IFM[72] Weight[75] Weight[74] Weight[73] Weight[72] N929 N928 N927 N926 N925 N924 N923 N922 CIM_DW_mult_uns_18
Xr828 IFM[71] IFM[70] IFM[69] IFM[68] Weight[71] Weight[70] Weight[69] Weight[68] N950 N949 N948 N947 N946 N945 N944 N943 CIM_DW_mult_uns_17
Xr830 IFM[67] IFM[66] IFM[65] IFM[64] Weight[67] Weight[66] Weight[65] Weight[64] N971 N970 N969 N968 N967 N966 N965 N964 CIM_DW_mult_uns_16
Xr832 IFM[63] IFM[62] IFM[61] IFM[60] Weight[63] Weight[62] Weight[61] Weight[60] N992 N991 N990 N989 N988 N987 N986 N985 CIM_DW_mult_uns_15
Xr834 IFM[59] IFM[58] IFM[57] IFM[56] Weight[59] Weight[58] Weight[57] Weight[56] N1013 N1012 N1011 N1010 N1009 N1008 N1007 N1006 CIM_DW_mult_uns_14
Xr836 IFM[55] IFM[54] IFM[53] IFM[52] Weight[55] Weight[54] Weight[53] Weight[52] N1034 N1033 N1032 N1031 N1030 N1029 N1028 N1027 CIM_DW_mult_uns_13
Xr838 IFM[51] IFM[50] IFM[49] IFM[48] Weight[51] Weight[50] Weight[49] Weight[48] N1055 N1054 N1053 N1052 N1051 N1050 N1049 N1048 CIM_DW_mult_uns_12
Xr840 IFM[47] IFM[46] IFM[45] IFM[44] Weight[47] Weight[46] Weight[45] Weight[44] N1076 N1075 N1074 N1073 N1072 N1071 N1070 N1069 CIM_DW_mult_uns_11
Xr842 IFM[43] IFM[42] IFM[41] IFM[40] Weight[43] Weight[42] Weight[41] Weight[40] N1097 N1096 N1095 N1094 N1093 N1092 N1091 N1090 CIM_DW_mult_uns_10
Xr844 IFM[39] IFM[38] IFM[37] IFM[36] Weight[39] Weight[38] Weight[37] Weight[36] N1118 N1117 N1116 N1115 N1114 N1113 N1112 N1111 CIM_DW_mult_uns_9
Xr846 IFM[35] IFM[34] IFM[33] IFM[32] Weight[35] Weight[34] Weight[33] Weight[32] N1139 N1138 N1137 N1136 N1135 N1134 N1133 N1132 CIM_DW_mult_uns_8
Xr848 IFM[31] IFM[30] IFM[29] IFM[28] Weight[31] Weight[30] Weight[29] Weight[28] N1160 N1159 N1158 N1157 N1156 N1155 N1154 N1153 CIM_DW_mult_uns_7
Xr850 IFM[27] IFM[26] IFM[25] IFM[24] Weight[27] Weight[26] Weight[25] Weight[24] N1181 N1180 N1179 N1178 N1177 N1176 N1175 N1174 CIM_DW_mult_uns_6
Xr852 IFM[23] IFM[22] IFM[21] IFM[20] Weight[23] Weight[22] Weight[21] Weight[20] N1202 N1201 N1200 N1199 N1198 N1197 N1196 N1195 CIM_DW_mult_uns_5
Xr854 IFM[19] IFM[18] IFM[17] IFM[16] Weight[19] Weight[18] Weight[17] Weight[16] N1223 N1222 N1221 N1220 N1219 N1218 N1217 N1216 CIM_DW_mult_uns_4
Xr856 IFM[15] IFM[14] IFM[13] IFM[12] Weight[15] Weight[14] Weight[13] Weight[12] N1244 N1243 N1242 N1241 N1240 N1239 N1238 N1237 CIM_DW_mult_uns_3
Xr858 IFM[11] IFM[10] IFM[9] IFM[8] Weight[11] Weight[10] Weight[9] Weight[8] N1265 N1264 N1263 N1262 N1261 N1260 N1259 N1258 CIM_DW_mult_uns_2
Xr860 IFM[7] IFM[6] IFM[5] IFM[4] Weight[7] Weight[6] Weight[5] Weight[4] N1286 N1285 N1284 N1283 N1282 N1281 N1280 N1279 CIM_DW_mult_uns_1
Xr862 IFM[3] IFM[2] IFM[1] IFM[0] Weight[3] Weight[2] Weight[1] Weight[0] N1307 N1306 N1305 N1304 N1303 N1302 N1301 N1300 CIM_DW_mult_uns_0
Xadd_2_root_r893 n1254 n1254 N1045 N1044 N1043 N1042 N1041 N1040 N1039 N1038 N1037 N1036 n1212 n1254 n1254 N1024 N1023 N1022 N1021 N1020 N1019 N1018 N1017 N1016 N1015 n1198 n1254 SYNOPSYS_UNCONNECTED_1 N1193 N1192 N1191 N1190 N1189 N1188 N1187 N1186 N1185 N1184 N1183 N1182 CIM_DW01_add_2
Xadd_1_root_r893 n1254 n1254 add_4_root_r893_SUM_10_ add_4_root_r893_SUM_9_ add_4_root_r893_SUM_8_ add_4_root_r893_SUM_7_ add_4_root_r893_SUM_6_ add_4_root_r893_SUM_5_ add_4_root_r893_SUM_4_ add_4_root_r893_SUM_3_ add_4_root_r893_SUM_2_ add_4_root_r893_SUM_1_ n1213 n1254 n1254 add_5_root_r893_SUM_10_ add_5_root_r893_SUM_9_ add_5_root_r893_SUM_8_ add_5_root_r893_SUM_7_ add_5_root_r893_SUM_6_ add_5_root_r893_SUM_5_ add_5_root_r893_SUM_4_ add_5_root_r893_SUM_3_ add_5_root_r893_SUM_2_ add_5_root_r893_SUM_1_ n1199 n1254 SYNOPSYS_UNCONNECTED_2 N1277 N1276 N1275 N1274 N1273 N1272 N1271 N1270 N1269 N1268 N1267 N1266 CIM_DW01_add_1
Xadd_0_root_r893 n1254 N1193 N1192 N1191 N1190 N1189 N1188 N1187 N1186 N1185 N1184 N1183 N1182 n1254 N1277 N1276 N1275 N1274 N1273 N1272 N1271 N1270 N1269 N1268 N1267 N1266 n1254 N1320 N1319 N1318 N1317 N1316 N1315 N1314 N1313 N1312 N1311 N1310 N1309 N1308 CIM_DW01_add_0
Xadd_6_root_r893_U1_1 N784 add_6_root_r893_B_1_ n1211 n1880 n1879 FAx1_ASAP7_75t_R
Xadd_6_root_r893_U1_2 N785 add_6_root_r893_B_2_ n1897 n1882 n1881 FAx1_ASAP7_75t_R
Xadd_6_root_r893_U1_3 N786 add_6_root_r893_B_3_ n1898 n1884 n1883 FAx1_ASAP7_75t_R
Xadd_6_root_r893_U1_4 N787 add_6_root_r893_B_4_ n1899 n1886 n1885 FAx1_ASAP7_75t_R
Xadd_6_root_r893_U1_5 N788 add_6_root_r893_B_5_ n1900 n1888 n1887 FAx1_ASAP7_75t_R
Xadd_6_root_r893_U1_6 N789 add_6_root_r893_B_6_ n1901 n1890 n1889 FAx1_ASAP7_75t_R
Xadd_6_root_r893_U1_7 N790 add_6_root_r893_B_7_ n1902 n1892 n1891 FAx1_ASAP7_75t_R
Xadd_6_root_r893_U1_8 N791 add_6_root_r893_B_8_ n1903 n1894 n1893 FAx1_ASAP7_75t_R
Xadd_6_root_r893_U1_9 N792 add_6_root_r893_B_9_ n1904 n1896 n1895 FAx1_ASAP7_75t_R
Xadd_3_root_r893_U1_1 N805 N763 n1210 n1854 n1853 FAx1_ASAP7_75t_R
Xadd_3_root_r893_U1_2 N806 N764 n1871 n1856 n1855 FAx1_ASAP7_75t_R
Xadd_3_root_r893_U1_3 N807 N765 n1872 n1858 n1857 FAx1_ASAP7_75t_R
Xadd_3_root_r893_U1_4 N808 N766 n1873 n1860 n1859 FAx1_ASAP7_75t_R
Xadd_3_root_r893_U1_5 N809 N767 n1874 n1862 n1861 FAx1_ASAP7_75t_R
Xadd_3_root_r893_U1_6 N810 N768 n1875 n1864 n1863 FAx1_ASAP7_75t_R
Xadd_3_root_r893_U1_7 N811 N769 n1876 n1866 n1865 FAx1_ASAP7_75t_R
Xadd_3_root_r893_U1_8 N812 N770 n1877 n1868 n1867 FAx1_ASAP7_75t_R
Xadd_3_root_r893_U1_9 N813 N771 n1878 n1870 n1869 FAx1_ASAP7_75t_R
Xadd_4_root_r893_U1_1 N1057 N1204 n1209 n1828 n1827 FAx1_ASAP7_75t_R
Xadd_4_root_r893_U1_2 N1058 N1205 n1845 n1830 n1829 FAx1_ASAP7_75t_R
Xadd_4_root_r893_U1_3 N1059 N1206 n1846 n1832 n1831 FAx1_ASAP7_75t_R
Xadd_4_root_r893_U1_4 N1060 N1207 n1847 n1834 n1833 FAx1_ASAP7_75t_R
Xadd_4_root_r893_U1_5 N1061 N1208 n1848 n1836 n1835 FAx1_ASAP7_75t_R
Xadd_4_root_r893_U1_6 N1062 N1209 n1849 n1838 n1837 FAx1_ASAP7_75t_R
Xadd_4_root_r893_U1_7 N1063 N1210 n1850 n1840 n1839 FAx1_ASAP7_75t_R
Xadd_4_root_r893_U1_8 N1064 N1211 n1851 n1842 n1841 FAx1_ASAP7_75t_R
Xadd_4_root_r893_U1_9 N1065 N1212 n1852 n1844 n1843 FAx1_ASAP7_75t_R
Xadd_9_root_r893_U1_1 N889 N868 n1207 n1805 n1804 FAx1_ASAP7_75t_R
Xadd_9_root_r893_U1_2 N890 N869 n1820 n1807 n1806 FAx1_ASAP7_75t_R
Xadd_9_root_r893_U1_3 N891 N870 n1821 n1809 n1808 FAx1_ASAP7_75t_R
Xadd_9_root_r893_U1_4 N892 N871 n1822 n1811 n1810 FAx1_ASAP7_75t_R
Xadd_9_root_r893_U1_5 N893 N872 n1823 n1813 n1812 FAx1_ASAP7_75t_R
Xadd_9_root_r893_U1_6 N894 N873 n1824 n1815 n1814 FAx1_ASAP7_75t_R
Xadd_9_root_r893_U1_7 N895 N874 n1825 n1817 n1816 FAx1_ASAP7_75t_R
Xadd_9_root_r893_U1_8 N896 N875 n1826 n1819 n1818 FAx1_ASAP7_75t_R
Xadd_10_root_r893_U1_1 N973 N847 n1206 n1782 n1781 FAx1_ASAP7_75t_R
Xadd_10_root_r893_U1_2 N974 N848 n1797 n1784 n1783 FAx1_ASAP7_75t_R
Xadd_10_root_r893_U1_3 N975 N849 n1798 n1786 n1785 FAx1_ASAP7_75t_R
Xadd_10_root_r893_U1_4 N976 N850 n1799 n1788 n1787 FAx1_ASAP7_75t_R
Xadd_10_root_r893_U1_5 N977 N851 n1800 n1790 n1789 FAx1_ASAP7_75t_R
Xadd_10_root_r893_U1_6 N978 N852 n1801 n1792 n1791 FAx1_ASAP7_75t_R
Xadd_10_root_r893_U1_7 N979 N853 n1802 n1794 n1793 FAx1_ASAP7_75t_R
Xadd_10_root_r893_U1_8 N980 N854 n1803 n1796 n1795 FAx1_ASAP7_75t_R
Xadd_29_root_r893_U1_1 N818 N986 n1241 n1762 n1761 FAx1_ASAP7_75t_R
Xadd_29_root_r893_U1_2 N819 N987 n1775 n1764 n1763 FAx1_ASAP7_75t_R
Xadd_29_root_r893_U1_3 N820 N988 n1776 n1766 n1765 FAx1_ASAP7_75t_R
Xadd_29_root_r893_U1_4 N821 N989 n1777 n1768 n1767 FAx1_ASAP7_75t_R
Xadd_29_root_r893_U1_5 N822 N990 n1778 n1770 n1769 FAx1_ASAP7_75t_R
Xadd_29_root_r893_U1_6 N823 N991 n1779 n1772 n1771 FAx1_ASAP7_75t_R
Xadd_29_root_r893_U1_7 N824 N992 n1780 n1774 n1773 FAx1_ASAP7_75t_R
Xadd_22_root_r893_U1_1 N19 N965 n1240 n1742 n1741 FAx1_ASAP7_75t_R
Xadd_22_root_r893_U1_2 N20 N966 n1755 n1744 n1743 FAx1_ASAP7_75t_R
Xadd_22_root_r893_U1_3 N21 N967 n1756 n1746 n1745 FAx1_ASAP7_75t_R
Xadd_22_root_r893_U1_4 N22 N968 n1757 n1748 n1747 FAx1_ASAP7_75t_R
Xadd_22_root_r893_U1_5 N23 N969 n1758 n1750 n1749 FAx1_ASAP7_75t_R
Xadd_22_root_r893_U1_6 N24 N970 n1759 n1752 n1751 FAx1_ASAP7_75t_R
Xadd_22_root_r893_U1_7 N25 N971 n1760 n1754 n1753 FAx1_ASAP7_75t_R
Xadd_20_root_r893_U1_1 N839 N1007 n1239 n1722 n1721 FAx1_ASAP7_75t_R
Xadd_20_root_r893_U1_2 N840 N1008 n1735 n1724 n1723 FAx1_ASAP7_75t_R
Xadd_20_root_r893_U1_3 N841 N1009 n1736 n1726 n1725 FAx1_ASAP7_75t_R
Xadd_20_root_r893_U1_4 N842 N1010 n1737 n1728 n1727 FAx1_ASAP7_75t_R
Xadd_20_root_r893_U1_5 N843 N1011 n1738 n1730 n1729 FAx1_ASAP7_75t_R
Xadd_20_root_r893_U1_6 N844 N1012 n1739 n1732 n1731 FAx1_ASAP7_75t_R
Xadd_20_root_r893_U1_7 N845 N1013 n1740 n1734 n1733 FAx1_ASAP7_75t_R
Xadd_19_root_r893_U1_1 N1049 N716 n1238 n1702 n1701 FAx1_ASAP7_75t_R
Xadd_19_root_r893_U1_2 N1050 N717 n1715 n1704 n1703 FAx1_ASAP7_75t_R
Xadd_19_root_r893_U1_3 N1051 N718 n1716 n1706 n1705 FAx1_ASAP7_75t_R
Xadd_19_root_r893_U1_4 N1052 N719 n1717 n1708 n1707 FAx1_ASAP7_75t_R
Xadd_19_root_r893_U1_5 N1053 N720 n1718 n1710 n1709 FAx1_ASAP7_75t_R
Xadd_19_root_r893_U1_6 N1054 N721 n1719 n1712 n1711 FAx1_ASAP7_75t_R
Xadd_19_root_r893_U1_7 N1055 N722 n1720 n1714 n1713 FAx1_ASAP7_75t_R
Xadd_14_root_r893_U1_1 N931 N826 n1205 n1679 n1678 FAx1_ASAP7_75t_R
Xadd_14_root_r893_U1_2 N932 N827 n1694 n1681 n1680 FAx1_ASAP7_75t_R
Xadd_14_root_r893_U1_3 N933 N828 n1695 n1683 n1682 FAx1_ASAP7_75t_R
Xadd_14_root_r893_U1_4 N934 N829 n1696 n1685 n1684 FAx1_ASAP7_75t_R
Xadd_14_root_r893_U1_5 N935 N830 n1697 n1687 n1686 FAx1_ASAP7_75t_R
Xadd_14_root_r893_U1_6 N936 N831 n1698 n1689 n1688 FAx1_ASAP7_75t_R
Xadd_14_root_r893_U1_7 N937 N832 n1699 n1691 n1690 FAx1_ASAP7_75t_R
Xadd_14_root_r893_U1_8 N938 N833 n1700 n1693 n1692 FAx1_ASAP7_75t_R
Xadd_15_root_r893_U1_1 N1175 N755 n1237 n1659 n1658 FAx1_ASAP7_75t_R
Xadd_15_root_r893_U1_2 N1176 N756 n1672 n1661 n1660 FAx1_ASAP7_75t_R
Xadd_15_root_r893_U1_3 N1177 N757 n1673 n1663 n1662 FAx1_ASAP7_75t_R
Xadd_15_root_r893_U1_4 N1178 N758 n1674 n1665 n1664 FAx1_ASAP7_75t_R
Xadd_15_root_r893_U1_5 N1179 N759 n1675 n1667 n1666 FAx1_ASAP7_75t_R
Xadd_15_root_r893_U1_6 N1180 N760 n1676 n1669 n1668 FAx1_ASAP7_75t_R
Xadd_15_root_r893_U1_7 N1181 N761 n1677 n1671 n1670 FAx1_ASAP7_75t_R
Xadd_26_root_r893_U1_1 N698 N902 n1236 n1639 n1638 FAx1_ASAP7_75t_R
Xadd_26_root_r893_U1_2 N699 N903 n1652 n1641 n1640 FAx1_ASAP7_75t_R
Xadd_26_root_r893_U1_3 N700 N904 n1653 n1643 n1642 FAx1_ASAP7_75t_R
Xadd_26_root_r893_U1_4 N701 N905 n1654 n1645 n1644 FAx1_ASAP7_75t_R
Xadd_26_root_r893_U1_5 N702 N906 n1655 n1647 n1646 FAx1_ASAP7_75t_R
Xadd_26_root_r893_U1_6 N703 N907 n1656 n1649 n1648 FAx1_ASAP7_75t_R
Xadd_26_root_r893_U1_7 N704 N908 n1657 n1651 n1650 FAx1_ASAP7_75t_R
Xadd_12_root_r893_U1_1 N1120 N1225 n1204 n1616 n1615 FAx1_ASAP7_75t_R
Xadd_12_root_r893_U1_2 N1121 N1226 n1631 n1618 n1617 FAx1_ASAP7_75t_R
Xadd_12_root_r893_U1_3 N1122 N1227 n1632 n1620 n1619 FAx1_ASAP7_75t_R
Xadd_12_root_r893_U1_4 N1123 N1228 n1633 n1622 n1621 FAx1_ASAP7_75t_R
Xadd_12_root_r893_U1_5 N1124 N1229 n1634 n1624 n1623 FAx1_ASAP7_75t_R
Xadd_12_root_r893_U1_6 N1125 N1230 n1635 n1626 n1625 FAx1_ASAP7_75t_R
Xadd_12_root_r893_U1_7 N1126 N1231 n1636 n1628 n1627 FAx1_ASAP7_75t_R
Xadd_12_root_r893_U1_8 N1127 N1232 n1637 n1630 n1629 FAx1_ASAP7_75t_R
Xadd_17_root_r893_U1_1 N1091 N1217 n1235 n1596 n1595 FAx1_ASAP7_75t_R
Xadd_17_root_r893_U1_2 N1092 N1218 n1609 n1598 n1597 FAx1_ASAP7_75t_R
Xadd_17_root_r893_U1_3 N1093 N1219 n1610 n1600 n1599 FAx1_ASAP7_75t_R
Xadd_17_root_r893_U1_4 N1094 N1220 n1611 n1602 n1601 FAx1_ASAP7_75t_R
Xadd_17_root_r893_U1_5 N1095 N1221 n1612 n1604 n1603 FAx1_ASAP7_75t_R
Xadd_17_root_r893_U1_6 N1096 N1222 n1613 n1606 n1605 FAx1_ASAP7_75t_R
Xadd_17_root_r893_U1_7 N1097 N1223 n1614 n1608 n1607 FAx1_ASAP7_75t_R
Xadd_21_root_r893_U1_1 N797 N1259 n1234 n1576 n1575 FAx1_ASAP7_75t_R
Xadd_21_root_r893_U1_2 N798 N1260 n1589 n1578 n1577 FAx1_ASAP7_75t_R
Xadd_21_root_r893_U1_3 N799 N1261 n1590 n1580 n1579 FAx1_ASAP7_75t_R
Xadd_21_root_r893_U1_4 N800 N1262 n1591 n1582 n1581 FAx1_ASAP7_75t_R
Xadd_21_root_r893_U1_5 N801 N1263 n1592 n1584 n1583 FAx1_ASAP7_75t_R
Xadd_21_root_r893_U1_6 N802 N1264 n1593 n1586 n1585 FAx1_ASAP7_75t_R
Xadd_21_root_r893_U1_7 N803 N1265 n1594 n1588 n1587 FAx1_ASAP7_75t_R
Xadd_11_root_r893_U1_1 N1246 N1099 n1203 n1553 n1552 FAx1_ASAP7_75t_R
Xadd_11_root_r893_U1_2 N1247 N1100 n1568 n1555 n1554 FAx1_ASAP7_75t_R
Xadd_11_root_r893_U1_3 N1248 N1101 n1569 n1557 n1556 FAx1_ASAP7_75t_R
Xadd_11_root_r893_U1_4 N1249 N1102 n1570 n1559 n1558 FAx1_ASAP7_75t_R
Xadd_11_root_r893_U1_5 N1250 N1103 n1571 n1561 n1560 FAx1_ASAP7_75t_R
Xadd_11_root_r893_U1_6 N1251 N1104 n1572 n1563 n1562 FAx1_ASAP7_75t_R
Xadd_11_root_r893_U1_7 N1252 N1105 n1573 n1565 n1564 FAx1_ASAP7_75t_R
Xadd_11_root_r893_U1_8 N1253 N1106 n1574 n1567 n1566 FAx1_ASAP7_75t_R
Xadd_18_root_r893_U1_1 N923 N1301 n1233 n1533 n1532 FAx1_ASAP7_75t_R
Xadd_18_root_r893_U1_2 N924 N1302 n1546 n1535 n1534 FAx1_ASAP7_75t_R
Xadd_18_root_r893_U1_3 N925 N1303 n1547 n1537 n1536 FAx1_ASAP7_75t_R
Xadd_18_root_r893_U1_4 N926 N1304 n1548 n1539 n1538 FAx1_ASAP7_75t_R
Xadd_18_root_r893_U1_5 N927 N1305 n1549 n1541 n1540 FAx1_ASAP7_75t_R
Xadd_18_root_r893_U1_6 N928 N1306 n1550 n1543 n1542 FAx1_ASAP7_75t_R
Xadd_18_root_r893_U1_7 N929 N1307 n1551 n1545 n1544 FAx1_ASAP7_75t_R
Xadd_24_root_r893_U1_1 N776 N1238 n1232 n1513 n1512 FAx1_ASAP7_75t_R
Xadd_24_root_r893_U1_2 N777 N1239 n1526 n1515 n1514 FAx1_ASAP7_75t_R
Xadd_24_root_r893_U1_3 N778 N1240 n1527 n1517 n1516 FAx1_ASAP7_75t_R
Xadd_24_root_r893_U1_4 N779 N1241 n1528 n1519 n1518 FAx1_ASAP7_75t_R
Xadd_24_root_r893_U1_5 N780 N1242 n1529 n1521 n1520 FAx1_ASAP7_75t_R
Xadd_24_root_r893_U1_6 N781 N1243 n1530 n1523 n1522 FAx1_ASAP7_75t_R
Xadd_24_root_r893_U1_7 N782 N1244 n1531 n1525 n1524 FAx1_ASAP7_75t_R
Xadd_7_root_r893_U1_1 N952 N1162 n1202 n1490 n1489 FAx1_ASAP7_75t_R
Xadd_7_root_r893_U1_2 N953 N1163 n1505 n1492 n1491 FAx1_ASAP7_75t_R
Xadd_7_root_r893_U1_3 N954 N1164 n1506 n1494 n1493 FAx1_ASAP7_75t_R
Xadd_7_root_r893_U1_4 N955 N1165 n1507 n1496 n1495 FAx1_ASAP7_75t_R
Xadd_7_root_r893_U1_5 N956 N1166 n1508 n1498 n1497 FAx1_ASAP7_75t_R
Xadd_7_root_r893_U1_6 N957 N1167 n1509 n1500 n1499 FAx1_ASAP7_75t_R
Xadd_7_root_r893_U1_7 N958 N1168 n1510 n1502 n1501 FAx1_ASAP7_75t_R
Xadd_7_root_r893_U1_8 N959 N1169 n1511 n1504 n1503 FAx1_ASAP7_75t_R
Xadd_28_root_r893_U1_1 N1028 N860 n1231 n1470 n1469 FAx1_ASAP7_75t_R
Xadd_28_root_r893_U1_2 N1029 N861 n1483 n1472 n1471 FAx1_ASAP7_75t_R
Xadd_28_root_r893_U1_3 N1030 N862 n1484 n1474 n1473 FAx1_ASAP7_75t_R
Xadd_28_root_r893_U1_4 N1031 N863 n1485 n1476 n1475 FAx1_ASAP7_75t_R
Xadd_28_root_r893_U1_5 N1032 N864 n1486 n1478 n1477 FAx1_ASAP7_75t_R
Xadd_28_root_r893_U1_6 N1033 N865 n1487 n1480 n1479 FAx1_ASAP7_75t_R
Xadd_28_root_r893_U1_7 N1034 N866 n1488 n1482 n1481 FAx1_ASAP7_75t_R
Xadd_27_root_r893_U1_1 N1070 N1112 n1230 n1450 n1449 FAx1_ASAP7_75t_R
Xadd_27_root_r893_U1_2 N1071 N1113 n1463 n1452 n1451 FAx1_ASAP7_75t_R
Xadd_27_root_r893_U1_3 N1072 N1114 n1464 n1454 n1453 FAx1_ASAP7_75t_R
Xadd_27_root_r893_U1_4 N1073 N1115 n1465 n1456 n1455 FAx1_ASAP7_75t_R
Xadd_27_root_r893_U1_5 N1074 N1116 n1466 n1458 n1457 FAx1_ASAP7_75t_R
Xadd_27_root_r893_U1_6 N1075 N1117 n1467 n1460 n1459 FAx1_ASAP7_75t_R
Xadd_27_root_r893_U1_7 N1076 N1118 n1468 n1462 n1461 FAx1_ASAP7_75t_R
Xadd_5_root_r893_U1_1 N1078 add_5_root_r893_B_1_ n1208 n1424 n1423 FAx1_ASAP7_75t_R
Xadd_5_root_r893_U1_2 N1079 add_5_root_r893_B_2_ n1441 n1426 n1425 FAx1_ASAP7_75t_R
Xadd_5_root_r893_U1_3 N1080 add_5_root_r893_B_3_ n1442 n1428 n1427 FAx1_ASAP7_75t_R
Xadd_5_root_r893_U1_4 N1081 add_5_root_r893_B_4_ n1443 n1430 n1429 FAx1_ASAP7_75t_R
Xadd_5_root_r893_U1_5 N1082 add_5_root_r893_B_5_ n1444 n1432 n1431 FAx1_ASAP7_75t_R
Xadd_5_root_r893_U1_6 N1083 add_5_root_r893_B_6_ n1445 n1434 n1433 FAx1_ASAP7_75t_R
Xadd_5_root_r893_U1_7 N1084 add_5_root_r893_B_7_ n1446 n1436 n1435 FAx1_ASAP7_75t_R
Xadd_5_root_r893_U1_8 N1085 add_5_root_r893_B_8_ n1447 n1438 n1437 FAx1_ASAP7_75t_R
Xadd_5_root_r893_U1_9 N1086 add_5_root_r893_B_9_ n1448 n1440 n1439 FAx1_ASAP7_75t_R
Xadd_8_root_r893_U1_1 N994 N910 n1201 n1401 n1400 FAx1_ASAP7_75t_R
Xadd_8_root_r893_U1_2 N995 N911 n1416 n1403 n1402 FAx1_ASAP7_75t_R
Xadd_8_root_r893_U1_3 N996 N912 n1417 n1405 n1404 FAx1_ASAP7_75t_R
Xadd_8_root_r893_U1_4 N997 N913 n1418 n1407 n1406 FAx1_ASAP7_75t_R
Xadd_8_root_r893_U1_5 N998 N914 n1419 n1409 n1408 FAx1_ASAP7_75t_R
Xadd_8_root_r893_U1_6 N999 N915 n1420 n1411 n1410 FAx1_ASAP7_75t_R
Xadd_8_root_r893_U1_7 N1000 N916 n1421 n1413 n1412 FAx1_ASAP7_75t_R
Xadd_8_root_r893_U1_8 N1001 N917 n1422 n1415 n1414 FAx1_ASAP7_75t_R
Xadd_23_root_r893_U1_1 N944 N1154 n1229 n1381 n1380 FAx1_ASAP7_75t_R
Xadd_23_root_r893_U1_2 N945 N1155 n1394 n1383 n1382 FAx1_ASAP7_75t_R
Xadd_23_root_r893_U1_3 N946 N1156 n1395 n1385 n1384 FAx1_ASAP7_75t_R
Xadd_23_root_r893_U1_4 N947 N1157 n1396 n1387 n1386 FAx1_ASAP7_75t_R
Xadd_23_root_r893_U1_5 N948 N1158 n1397 n1389 n1388 FAx1_ASAP7_75t_R
Xadd_23_root_r893_U1_6 N949 N1159 n1398 n1391 n1390 FAx1_ASAP7_75t_R
Xadd_23_root_r893_U1_7 N950 N1160 n1399 n1393 n1392 FAx1_ASAP7_75t_R
Xadd_30_root_r893_U1_1 N11 N735 n1228 n1361 n1360 FAx1_ASAP7_75t_R
Xadd_30_root_r893_U1_2 N12 N736 n1374 n1363 n1362 FAx1_ASAP7_75t_R
Xadd_30_root_r893_U1_3 N13 N737 n1375 n1365 n1364 FAx1_ASAP7_75t_R
Xadd_30_root_r893_U1_4 N14 N738 n1376 n1367 n1366 FAx1_ASAP7_75t_R
Xadd_30_root_r893_U1_5 N15 N739 n1377 n1369 n1368 FAx1_ASAP7_75t_R
Xadd_30_root_r893_U1_6 N16 N740 n1378 n1371 n1370 FAx1_ASAP7_75t_R
Xadd_30_root_r893_U1_7 N17 N741 n1379 n1373 n1372 FAx1_ASAP7_75t_R
Xadd_13_root_r893_U1_1 N1141 N1288 n1200 n1338 n1337 FAx1_ASAP7_75t_R
Xadd_13_root_r893_U1_2 N1142 N1289 n1353 n1340 n1339 FAx1_ASAP7_75t_R
Xadd_13_root_r893_U1_3 N1143 N1290 n1354 n1342 n1341 FAx1_ASAP7_75t_R
Xadd_13_root_r893_U1_4 N1144 N1291 n1355 n1344 n1343 FAx1_ASAP7_75t_R
Xadd_13_root_r893_U1_5 N1145 N1292 n1356 n1346 n1345 FAx1_ASAP7_75t_R
Xadd_13_root_r893_U1_6 N1146 N1293 n1357 n1348 n1347 FAx1_ASAP7_75t_R
Xadd_13_root_r893_U1_7 N1147 N1294 n1358 n1350 n1349 FAx1_ASAP7_75t_R
Xadd_13_root_r893_U1_8 N1148 N1295 n1359 n1352 n1351 FAx1_ASAP7_75t_R
Xadd_16_root_r893_U1_1 N881 N1133 n1227 n1318 n1317 FAx1_ASAP7_75t_R
Xadd_16_root_r893_U1_2 N882 N1134 n1331 n1320 n1319 FAx1_ASAP7_75t_R
Xadd_16_root_r893_U1_3 N883 N1135 n1332 n1322 n1321 FAx1_ASAP7_75t_R
Xadd_16_root_r893_U1_4 N884 N1136 n1333 n1324 n1323 FAx1_ASAP7_75t_R
Xadd_16_root_r893_U1_5 N885 N1137 n1334 n1326 n1325 FAx1_ASAP7_75t_R
Xadd_16_root_r893_U1_6 N886 N1138 n1335 n1328 n1327 FAx1_ASAP7_75t_R
Xadd_16_root_r893_U1_7 N887 N1139 n1336 n1330 n1329 FAx1_ASAP7_75t_R
Xadd_25_root_r893_U1_1 N1196 N1280 n1226 n1298 n1297 FAx1_ASAP7_75t_R
Xadd_25_root_r893_U1_2 N1197 N1281 n1311 n1300 n1299 FAx1_ASAP7_75t_R
Xadd_25_root_r893_U1_3 N1198 N1282 n1312 n1302 n1301 FAx1_ASAP7_75t_R
Xadd_25_root_r893_U1_4 N1199 N1283 n1313 n1304 n1303 FAx1_ASAP7_75t_R
Xadd_25_root_r893_U1_5 N1200 N1284 n1314 n1306 n1305 FAx1_ASAP7_75t_R
Xadd_25_root_r893_U1_6 N1201 N1285 n1315 n1308 n1307 FAx1_ASAP7_75t_R
Xadd_25_root_r893_U1_7 N1202 N1286 n1316 n1310 n1309 FAx1_ASAP7_75t_R
Xclk22_reg clk22 clk n1254 n1905 clk22 ASYNC_DFFHx1_ASAP7_75t_R
Xout_valid_reg n1906 clk n1905 n1254 out_valid ASYNC_DFFHx1_ASAP7_75t_R
Xstate_cs_reg n1261 clk n1905 n1254 state_cs ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_2__3_ n927 clk n1905 n1254 Weight[123] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_2__0_ n921 clk n1905 n1254 Weight[120] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_1__3_ n935 clk n1905 n1254 Weight[127] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_1__0_ n929 clk n1905 n1254 Weight[124] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_2__1_ n923 clk n1905 n1254 Weight[121] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_1__1_ n931 clk n1905 n1254 Weight[125] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_2__2_ n925 clk n1905 n1254 Weight[122] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_1__2_ n933 clk n1905 n1254 Weight[126] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_2__3_ n1183 clk n1905 n1254 IFM[123] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_2__2_ n1181 clk n1905 n1254 IFM[122] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_2__1_ n1179 clk n1905 n1254 IFM[121] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_2__0_ n1177 clk n1905 n1254 IFM[120] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_1__3_ n1191 clk n1905 n1254 IFM[127] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_1__2_ n1189 clk n1905 n1254 IFM[126] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_1__1_ n1187 clk n1905 n1254 IFM[125] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_1__0_ n1185 clk n1905 n1254 IFM[124] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_32__3_ n687 clk n1905 n1254 Weight[3] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_32__0_ n681 clk n1905 n1254 Weight[0] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_31__3_ n695 clk n1905 n1254 Weight[7] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_31__0_ n689 clk n1905 n1254 Weight[4] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_30__3_ n703 clk n1905 n1254 Weight[11] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_30__0_ n697 clk n1905 n1254 Weight[8] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_29__3_ n711 clk n1905 n1254 Weight[15] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_29__0_ n705 clk n1905 n1254 Weight[12] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_28__3_ n719 clk n1905 n1254 Weight[19] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_28__0_ n713 clk n1905 n1254 Weight[16] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_27__3_ n727 clk n1905 n1254 Weight[23] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_27__0_ n721 clk n1905 n1254 Weight[20] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_26__3_ n735 clk n1905 n1254 Weight[27] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_26__0_ n729 clk n1905 n1254 Weight[24] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_25__3_ n743 clk n1905 n1254 Weight[31] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_25__0_ n737 clk n1905 n1254 Weight[28] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_24__3_ n751 clk n1905 n1254 Weight[35] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_24__0_ n745 clk n1905 n1254 Weight[32] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_23__3_ n759 clk n1905 n1254 Weight[39] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_23__0_ n753 clk n1905 n1254 Weight[36] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_22__3_ n767 clk n1905 n1254 Weight[43] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_22__0_ n761 clk n1905 n1254 Weight[40] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_21__3_ n775 clk n1905 n1254 Weight[47] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_21__0_ n769 clk n1905 n1254 Weight[44] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_20__3_ n783 clk n1905 n1254 Weight[51] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_20__0_ n777 clk n1905 n1254 Weight[48] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_19__3_ n791 clk n1905 n1254 Weight[55] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_19__0_ n785 clk n1905 n1254 Weight[52] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_18__3_ n799 clk n1905 n1254 Weight[59] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_18__0_ n793 clk n1905 n1254 Weight[56] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_17__3_ n807 clk n1905 n1254 Weight[63] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_17__0_ n801 clk n1905 n1254 Weight[60] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_16__3_ n815 clk n1905 n1254 Weight[67] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_16__0_ n809 clk n1905 n1254 Weight[64] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_15__3_ n823 clk n1905 n1254 Weight[71] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_15__0_ n817 clk n1905 n1254 Weight[68] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_14__3_ n831 clk n1905 n1254 Weight[75] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_14__0_ n825 clk n1905 n1254 Weight[72] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_13__3_ n839 clk n1905 n1254 Weight[79] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_13__0_ n833 clk n1905 n1254 Weight[76] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_12__3_ n847 clk n1905 n1254 Weight[83] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_12__0_ n841 clk n1905 n1254 Weight[80] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_11__3_ n855 clk n1905 n1254 Weight[87] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_11__0_ n849 clk n1905 n1254 Weight[84] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_10__3_ n863 clk n1905 n1254 Weight[91] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_10__0_ n857 clk n1905 n1254 Weight[88] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_9__3_ n871 clk n1905 n1254 Weight[95] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_9__0_ n865 clk n1905 n1254 Weight[92] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_8__3_ n879 clk n1905 n1254 Weight[99] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_8__0_ n873 clk n1905 n1254 Weight[96] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_7__3_ n887 clk n1905 n1254 Weight[103] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_7__0_ n881 clk n1905 n1254 Weight[100] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_6__3_ n895 clk n1905 n1254 Weight[107] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_6__0_ n889 clk n1905 n1254 Weight[104] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_5__3_ n903 clk n1905 n1254 Weight[111] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_5__0_ n897 clk n1905 n1254 Weight[108] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_4__3_ n911 clk n1905 n1254 Weight[115] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_4__0_ n905 clk n1905 n1254 Weight[112] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_3__3_ n919 clk n1905 n1254 Weight[119] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_3__0_ n913 clk n1905 n1254 Weight[116] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_32__1_ n683 clk n1905 n1254 Weight[1] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_31__1_ n691 clk n1905 n1254 Weight[5] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_30__1_ n699 clk n1905 n1254 Weight[9] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_29__1_ n707 clk n1905 n1254 Weight[13] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_28__1_ n715 clk n1905 n1254 Weight[17] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_27__1_ n723 clk n1905 n1254 Weight[21] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_26__1_ n731 clk n1905 n1254 Weight[25] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_25__1_ n739 clk n1905 n1254 Weight[29] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_24__1_ n747 clk n1905 n1254 Weight[33] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_23__1_ n755 clk n1905 n1254 Weight[37] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_22__1_ n763 clk n1905 n1254 Weight[41] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_21__1_ n771 clk n1905 n1254 Weight[45] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_20__1_ n779 clk n1905 n1254 Weight[49] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_19__1_ n787 clk n1905 n1254 Weight[53] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_18__1_ n795 clk n1905 n1254 Weight[57] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_17__1_ n803 clk n1905 n1254 Weight[61] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_16__1_ n811 clk n1905 n1254 Weight[65] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_15__1_ n819 clk n1905 n1254 Weight[69] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_14__1_ n827 clk n1905 n1254 Weight[73] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_13__1_ n835 clk n1905 n1254 Weight[77] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_12__1_ n843 clk n1905 n1254 Weight[81] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_11__1_ n851 clk n1905 n1254 Weight[85] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_10__1_ n859 clk n1905 n1254 Weight[89] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_9__1_ n867 clk n1905 n1254 Weight[93] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_8__1_ n875 clk n1905 n1254 Weight[97] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_7__1_ n883 clk n1905 n1254 Weight[101] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_6__1_ n891 clk n1905 n1254 Weight[105] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_5__1_ n899 clk n1905 n1254 Weight[109] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_4__1_ n907 clk n1905 n1254 Weight[113] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_3__1_ n915 clk n1905 n1254 Weight[117] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_32__2_ n685 clk n1905 n1254 Weight[2] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_31__2_ n693 clk n1905 n1254 Weight[6] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_30__2_ n701 clk n1905 n1254 Weight[10] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_29__2_ n709 clk n1905 n1254 Weight[14] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_28__2_ n717 clk n1905 n1254 Weight[18] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_27__2_ n725 clk n1905 n1254 Weight[22] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_26__2_ n733 clk n1905 n1254 Weight[26] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_25__2_ n741 clk n1905 n1254 Weight[30] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_24__2_ n749 clk n1905 n1254 Weight[34] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_23__2_ n757 clk n1905 n1254 Weight[38] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_22__2_ n765 clk n1905 n1254 Weight[42] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_21__2_ n773 clk n1905 n1254 Weight[46] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_20__2_ n781 clk n1905 n1254 Weight[50] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_19__2_ n789 clk n1905 n1254 Weight[54] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_18__2_ n797 clk n1905 n1254 Weight[58] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_17__2_ n805 clk n1905 n1254 Weight[62] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_16__2_ n813 clk n1905 n1254 Weight[66] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_15__2_ n821 clk n1905 n1254 Weight[70] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_14__2_ n829 clk n1905 n1254 Weight[74] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_13__2_ n837 clk n1905 n1254 Weight[78] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_12__2_ n845 clk n1905 n1254 Weight[82] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_11__2_ n853 clk n1905 n1254 Weight[86] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_10__2_ n861 clk n1905 n1254 Weight[90] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_9__2_ n869 clk n1905 n1254 Weight[94] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_8__2_ n877 clk n1905 n1254 Weight[98] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_7__2_ n885 clk n1905 n1254 Weight[102] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_6__2_ n893 clk n1905 n1254 Weight[106] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_5__2_ n901 clk n1905 n1254 Weight[110] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_4__2_ n909 clk n1905 n1254 Weight[114] ASYNC_DFFHx1_ASAP7_75t_R
XWeight_reg_3__2_ n917 clk n1905 n1254 Weight[118] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_32__3_ n943 clk n1905 n1254 IFM[3] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_32__2_ n941 clk n1905 n1254 IFM[2] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_32__1_ n939 clk n1905 n1254 IFM[1] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_32__0_ n937 clk n1905 n1254 IFM[0] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_31__3_ n951 clk n1905 n1254 IFM[7] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_31__2_ n949 clk n1905 n1254 IFM[6] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_31__1_ n947 clk n1905 n1254 IFM[5] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_31__0_ n945 clk n1905 n1254 IFM[4] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_30__3_ n959 clk n1905 n1254 IFM[11] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_30__2_ n957 clk n1905 n1254 IFM[10] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_30__1_ n955 clk n1905 n1254 IFM[9] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_30__0_ n953 clk n1905 n1254 IFM[8] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_29__3_ n967 clk n1905 n1254 IFM[15] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_29__2_ n965 clk n1905 n1254 IFM[14] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_29__1_ n963 clk n1905 n1254 IFM[13] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_29__0_ n961 clk n1905 n1254 IFM[12] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_28__3_ n975 clk n1905 n1254 IFM[19] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_28__2_ n973 clk n1905 n1254 IFM[18] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_28__1_ n971 clk n1905 n1254 IFM[17] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_28__0_ n969 clk n1905 n1254 IFM[16] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_27__3_ n983 clk n1905 n1254 IFM[23] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_27__2_ n981 clk n1905 n1254 IFM[22] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_27__1_ n979 clk n1905 n1254 IFM[21] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_27__0_ n977 clk n1905 n1254 IFM[20] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_26__3_ n991 clk n1905 n1254 IFM[27] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_26__2_ n989 clk n1905 n1254 IFM[26] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_26__1_ n987 clk n1905 n1254 IFM[25] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_26__0_ n985 clk n1905 n1254 IFM[24] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_25__3_ n999 clk n1905 n1254 IFM[31] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_25__2_ n997 clk n1905 n1254 IFM[30] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_25__1_ n995 clk n1905 n1254 IFM[29] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_25__0_ n993 clk n1905 n1254 IFM[28] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_24__3_ n1007 clk n1905 n1254 IFM[35] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_24__2_ n1005 clk n1905 n1254 IFM[34] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_24__1_ n1003 clk n1905 n1254 IFM[33] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_24__0_ n1001 clk n1905 n1254 IFM[32] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_23__3_ n1015 clk n1905 n1254 IFM[39] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_23__2_ n1013 clk n1905 n1254 IFM[38] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_23__1_ n1011 clk n1905 n1254 IFM[37] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_23__0_ n1009 clk n1905 n1254 IFM[36] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_22__3_ n1023 clk n1905 n1254 IFM[43] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_22__2_ n1021 clk n1905 n1254 IFM[42] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_22__1_ n1019 clk n1905 n1254 IFM[41] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_22__0_ n1017 clk n1905 n1254 IFM[40] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_21__3_ n1031 clk n1905 n1254 IFM[47] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_21__2_ n1029 clk n1905 n1254 IFM[46] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_21__1_ n1027 clk n1905 n1254 IFM[45] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_21__0_ n1025 clk n1905 n1254 IFM[44] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_20__3_ n1039 clk n1905 n1254 IFM[51] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_20__2_ n1037 clk n1905 n1254 IFM[50] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_20__1_ n1035 clk n1905 n1254 IFM[49] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_20__0_ n1033 clk n1905 n1254 IFM[48] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_19__3_ n1047 clk n1905 n1254 IFM[55] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_19__2_ n1045 clk n1905 n1254 IFM[54] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_19__1_ n1043 clk n1905 n1254 IFM[53] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_19__0_ n1041 clk n1905 n1254 IFM[52] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_18__3_ n1055 clk n1905 n1254 IFM[59] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_18__2_ n1053 clk n1905 n1254 IFM[58] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_18__1_ n1051 clk n1905 n1254 IFM[57] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_18__0_ n1049 clk n1905 n1254 IFM[56] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_17__3_ n1063 clk n1905 n1254 IFM[63] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_17__2_ n1061 clk n1905 n1254 IFM[62] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_17__1_ n1059 clk n1905 n1254 IFM[61] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_17__0_ n1057 clk n1905 n1254 IFM[60] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_16__3_ n1071 clk n1905 n1254 IFM[67] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_16__2_ n1069 clk n1905 n1254 IFM[66] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_16__1_ n1067 clk n1905 n1254 IFM[65] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_16__0_ n1065 clk n1905 n1254 IFM[64] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_15__3_ n1079 clk n1905 n1254 IFM[71] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_15__2_ n1077 clk n1905 n1254 IFM[70] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_15__1_ n1075 clk n1905 n1254 IFM[69] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_15__0_ n1073 clk n1905 n1254 IFM[68] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_14__3_ n1087 clk n1905 n1254 IFM[75] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_14__2_ n1085 clk n1905 n1254 IFM[74] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_14__1_ n1083 clk n1905 n1254 IFM[73] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_14__0_ n1081 clk n1905 n1254 IFM[72] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_13__3_ n1095 clk n1905 n1254 IFM[79] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_13__2_ n1093 clk n1905 n1254 IFM[78] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_13__1_ n1091 clk n1905 n1254 IFM[77] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_13__0_ n1089 clk n1905 n1254 IFM[76] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_12__3_ n1103 clk n1905 n1254 IFM[83] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_12__2_ n1101 clk n1905 n1254 IFM[82] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_12__1_ n1099 clk n1905 n1254 IFM[81] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_12__0_ n1097 clk n1905 n1254 IFM[80] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_11__3_ n1111 clk n1905 n1254 IFM[87] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_11__2_ n1109 clk n1905 n1254 IFM[86] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_11__1_ n1107 clk n1905 n1254 IFM[85] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_11__0_ n1105 clk n1905 n1254 IFM[84] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_10__3_ n1119 clk n1905 n1254 IFM[91] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_10__2_ n1117 clk n1905 n1254 IFM[90] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_10__1_ n1115 clk n1905 n1254 IFM[89] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_10__0_ n1113 clk n1905 n1254 IFM[88] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_9__3_ n1127 clk n1905 n1254 IFM[95] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_9__2_ n1125 clk n1905 n1254 IFM[94] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_9__1_ n1123 clk n1905 n1254 IFM[93] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_9__0_ n1121 clk n1905 n1254 IFM[92] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_8__3_ n1135 clk n1905 n1254 IFM[99] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_8__2_ n1133 clk n1905 n1254 IFM[98] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_8__1_ n1131 clk n1905 n1254 IFM[97] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_8__0_ n1129 clk n1905 n1254 IFM[96] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_7__3_ n1143 clk n1905 n1254 IFM[103] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_7__2_ n1141 clk n1905 n1254 IFM[102] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_7__1_ n1139 clk n1905 n1254 IFM[101] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_7__0_ n1137 clk n1905 n1254 IFM[100] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_6__3_ n1151 clk n1905 n1254 IFM[107] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_6__2_ n1149 clk n1905 n1254 IFM[106] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_6__1_ n1147 clk n1905 n1254 IFM[105] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_6__0_ n1145 clk n1905 n1254 IFM[104] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_5__3_ n1159 clk n1905 n1254 IFM[111] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_5__2_ n1157 clk n1905 n1254 IFM[110] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_5__1_ n1155 clk n1905 n1254 IFM[109] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_5__0_ n1153 clk n1905 n1254 IFM[108] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_4__3_ n1167 clk n1905 n1254 IFM[115] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_4__2_ n1165 clk n1905 n1254 IFM[114] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_4__1_ n1163 clk n1905 n1254 IFM[113] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_4__0_ n1161 clk n1905 n1254 IFM[112] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_3__3_ n1175 clk n1905 n1254 IFM[119] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_3__2_ n1173 clk n1905 n1254 IFM[118] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_3__1_ n1171 clk n1905 n1254 IFM[117] ASYNC_DFFHx1_ASAP7_75t_R
XIFM_reg_3__0_ n1169 clk n1905 n1254 IFM[116] ASYNC_DFFHx1_ASAP7_75t_R
XU1089 n1254 TIELOx1_ASAP7_75t_R
XU1090 n1224 n1252 n1198 XOR2xp5_ASAP7_75t_R
XU1091 n1222 n1250 n1199 XOR2xp5_ASAP7_75t_R
XU1092 n1218 n1243 n1200 AND2x2_ASAP7_75t_R
XU1093 n1214 n1242 n1201 AND2x2_ASAP7_75t_R
XU1094 n1217 n1248 n1202 AND2x2_ASAP7_75t_R
XU1095 n1216 n1246 n1203 AND2x2_ASAP7_75t_R
XU1096 n1221 n1249 n1204 AND2x2_ASAP7_75t_R
XU1097 n1220 n1247 n1205 AND2x2_ASAP7_75t_R
XU1098 n1219 n1245 n1206 AND2x2_ASAP7_75t_R
XU1099 n1215 n1244 n1207 AND2x2_ASAP7_75t_R
XU1100 n1222 n1250 n1208 AND2x2_ASAP7_75t_R
XU1101 n1223 n1251 n1209 AND2x2_ASAP7_75t_R
XU1102 n1224 n1252 n1210 AND2x2_ASAP7_75t_R
XU1103 n1225 n1253 n1211 AND2x2_ASAP7_75t_R
XU1104 n1225 n1253 n1212 XOR2xp5_ASAP7_75t_R
XU1105 n1223 n1251 n1213 XOR2xp5_ASAP7_75t_R
XU1106 N10 N734 n1214 XOR2xp5_ASAP7_75t_R
XU1107 N18 N964 n1215 XOR2xp5_ASAP7_75t_R
XU1108 N775 N1237 n1216 XOR2xp5_ASAP7_75t_R
XU1109 N1069 N1111 n1217 XOR2xp5_ASAP7_75t_R
XU1110 N1195 N1279 n1218 XOR2xp5_ASAP7_75t_R
XU1111 N817 N985 n1219 XOR2xp5_ASAP7_75t_R
XU1112 N697 N901 n1220 XOR2xp5_ASAP7_75t_R
XU1113 N796 N1258 n1221 XOR2xp5_ASAP7_75t_R
XU1114 n1218 n1243 n1222 XOR2xp5_ASAP7_75t_R
XU1115 n1219 n1245 n1223 XOR2xp5_ASAP7_75t_R
XU1116 n1220 n1247 n1224 XOR2xp5_ASAP7_75t_R
XU1117 n1221 n1249 n1225 XOR2xp5_ASAP7_75t_R
XU1118 N1195 N1279 n1226 AND2x2_ASAP7_75t_R
XU1119 N880 N1132 n1227 AND2x2_ASAP7_75t_R
XU1120 N10 N734 n1228 AND2x2_ASAP7_75t_R
XU1121 N943 N1153 n1229 AND2x2_ASAP7_75t_R
XU1122 N1069 N1111 n1230 AND2x2_ASAP7_75t_R
XU1123 N1027 N859 n1231 AND2x2_ASAP7_75t_R
XU1124 N775 N1237 n1232 AND2x2_ASAP7_75t_R
XU1125 N922 N1300 n1233 AND2x2_ASAP7_75t_R
XU1126 N796 N1258 n1234 AND2x2_ASAP7_75t_R
XU1127 N1090 N1216 n1235 AND2x2_ASAP7_75t_R
XU1128 N697 N901 n1236 AND2x2_ASAP7_75t_R
XU1129 N1174 N754 n1237 AND2x2_ASAP7_75t_R
XU1130 N1048 N715 n1238 AND2x2_ASAP7_75t_R
XU1131 N838 N1006 n1239 AND2x2_ASAP7_75t_R
XU1132 N18 N964 n1240 AND2x2_ASAP7_75t_R
XU1133 N817 N985 n1241 AND2x2_ASAP7_75t_R
XU1134 N943 N1153 n1242 XOR2xp5_ASAP7_75t_R
XU1135 N880 N1132 n1243 XOR2xp5_ASAP7_75t_R
XU1136 N838 N1006 n1244 XOR2xp5_ASAP7_75t_R
XU1137 N1048 N715 n1245 XOR2xp5_ASAP7_75t_R
XU1138 N922 N1300 n1246 XOR2xp5_ASAP7_75t_R
XU1139 N1174 N754 n1247 XOR2xp5_ASAP7_75t_R
XU1140 N1027 N859 n1248 XOR2xp5_ASAP7_75t_R
XU1141 N1090 N1216 n1249 XOR2xp5_ASAP7_75t_R
XU1142 n1214 n1242 n1250 XOR2xp5_ASAP7_75t_R
XU1143 n1215 n1244 n1251 XOR2xp5_ASAP7_75t_R
XU1144 n1216 n1246 n1252 XOR2xp5_ASAP7_75t_R
XU1145 n1217 n1248 n1253 XOR2xp5_ASAP7_75t_R
XU1146 rst_n n1905 INVx6_ASAP7_75t_R
XU1147 weight_valid n1255 INVx1_ASAP7_75t_R
XU1148 weight_valid n1256 INVx1_ASAP7_75t_R
XU1149 weight_valid n1257 INVx1_ASAP7_75t_R
XU1150 weight_valid n1258 INVx1_ASAP7_75t_R
XU1151 weight_valid n1259 INVx1_ASAP7_75t_R
XU1152 weight_valid n1260 INVx1_ASAP7_75t_R
XU1153 weight_valid Weight[0] n126 NOR2xp33_ASAP7_75t_R
XU1154 In_Weight[127] n1255 n125 NOR2xp33_ASAP7_75t_R
XU1155 weight_valid Weight[1] n129 NOR2xp33_ASAP7_75t_R
XU1156 In_Weight[126] n1255 n128 NOR2xp33_ASAP7_75t_R
XU1157 weight_valid Weight[2] n131 NOR2xp33_ASAP7_75t_R
XU1158 In_Weight[125] n1255 n130 NOR2xp33_ASAP7_75t_R
XU1159 weight_valid Weight[3] n133 NOR2xp33_ASAP7_75t_R
XU1160 In_Weight[124] n1255 n132 NOR2xp33_ASAP7_75t_R
XU1161 weight_valid Weight[4] n135 NOR2xp33_ASAP7_75t_R
XU1162 In_Weight[123] n1255 n134 NOR2xp33_ASAP7_75t_R
XU1163 weight_valid Weight[5] n137 NOR2xp33_ASAP7_75t_R
XU1164 In_Weight[122] n1255 n136 NOR2xp33_ASAP7_75t_R
XU1165 weight_valid Weight[6] n139 NOR2xp33_ASAP7_75t_R
XU1166 In_Weight[121] n1255 n138 NOR2xp33_ASAP7_75t_R
XU1167 weight_valid Weight[7] n141 NOR2xp33_ASAP7_75t_R
XU1168 In_Weight[120] n1255 n140 NOR2xp33_ASAP7_75t_R
XU1169 weight_valid Weight[8] n143 NOR2xp33_ASAP7_75t_R
XU1170 In_Weight[119] n1255 n142 NOR2xp33_ASAP7_75t_R
XU1171 weight_valid Weight[9] n145 NOR2xp33_ASAP7_75t_R
XU1172 In_Weight[118] n1255 n144 NOR2xp33_ASAP7_75t_R
XU1173 weight_valid Weight[10] n147 NOR2xp33_ASAP7_75t_R
XU1174 In_Weight[117] n1255 n146 NOR2xp33_ASAP7_75t_R
XU1175 weight_valid Weight[11] n149 NOR2xp33_ASAP7_75t_R
XU1176 In_Weight[116] n1255 n148 NOR2xp33_ASAP7_75t_R
XU1177 weight_valid Weight[12] n151 NOR2xp33_ASAP7_75t_R
XU1178 In_Weight[115] n1256 n150 NOR2xp33_ASAP7_75t_R
XU1179 weight_valid Weight[13] n153 NOR2xp33_ASAP7_75t_R
XU1180 In_Weight[114] n1256 n152 NOR2xp33_ASAP7_75t_R
XU1181 weight_valid Weight[14] n155 NOR2xp33_ASAP7_75t_R
XU1182 In_Weight[113] n1256 n154 NOR2xp33_ASAP7_75t_R
XU1183 weight_valid Weight[15] n157 NOR2xp33_ASAP7_75t_R
XU1184 In_Weight[112] n1256 n156 NOR2xp33_ASAP7_75t_R
XU1185 weight_valid Weight[16] n159 NOR2xp33_ASAP7_75t_R
XU1186 In_Weight[111] n1256 n158 NOR2xp33_ASAP7_75t_R
XU1187 weight_valid Weight[17] n161 NOR2xp33_ASAP7_75t_R
XU1188 In_Weight[110] n1256 n160 NOR2xp33_ASAP7_75t_R
XU1189 weight_valid Weight[18] n163 NOR2xp33_ASAP7_75t_R
XU1190 In_Weight[109] n1256 n162 NOR2xp33_ASAP7_75t_R
XU1191 weight_valid Weight[19] n165 NOR2xp33_ASAP7_75t_R
XU1192 In_Weight[108] n1256 n164 NOR2xp33_ASAP7_75t_R
XU1193 weight_valid Weight[20] n167 NOR2xp33_ASAP7_75t_R
XU1194 In_Weight[107] n1256 n166 NOR2xp33_ASAP7_75t_R
XU1195 weight_valid Weight[21] n169 NOR2xp33_ASAP7_75t_R
XU1196 In_Weight[106] n1256 n168 NOR2xp33_ASAP7_75t_R
XU1197 weight_valid Weight[22] n171 NOR2xp33_ASAP7_75t_R
XU1198 In_Weight[105] n1256 n170 NOR2xp33_ASAP7_75t_R
XU1199 weight_valid Weight[23] n173 NOR2xp33_ASAP7_75t_R
XU1200 In_Weight[104] n1256 n172 NOR2xp33_ASAP7_75t_R
XU1201 weight_valid Weight[24] n175 NOR2xp33_ASAP7_75t_R
XU1202 In_Weight[103] n1257 n174 NOR2xp33_ASAP7_75t_R
XU1203 weight_valid Weight[25] n177 NOR2xp33_ASAP7_75t_R
XU1204 In_Weight[102] n1257 n176 NOR2xp33_ASAP7_75t_R
XU1205 weight_valid Weight[26] n179 NOR2xp33_ASAP7_75t_R
XU1206 In_Weight[101] n1257 n178 NOR2xp33_ASAP7_75t_R
XU1207 weight_valid Weight[27] n181 NOR2xp33_ASAP7_75t_R
XU1208 In_Weight[100] n1257 n180 NOR2xp33_ASAP7_75t_R
XU1209 weight_valid Weight[28] n183 NOR2xp33_ASAP7_75t_R
XU1210 In_Weight[99] n1257 n182 NOR2xp33_ASAP7_75t_R
XU1211 weight_valid Weight[29] n185 NOR2xp33_ASAP7_75t_R
XU1212 In_Weight[98] n1257 n184 NOR2xp33_ASAP7_75t_R
XU1213 weight_valid Weight[30] n187 NOR2xp33_ASAP7_75t_R
XU1214 In_Weight[97] n1257 n186 NOR2xp33_ASAP7_75t_R
XU1215 weight_valid Weight[31] n189 NOR2xp33_ASAP7_75t_R
XU1216 In_Weight[96] n1257 n188 NOR2xp33_ASAP7_75t_R
XU1217 weight_valid Weight[32] n191 NOR2xp33_ASAP7_75t_R
XU1218 In_Weight[95] n1257 n190 NOR2xp33_ASAP7_75t_R
XU1219 weight_valid Weight[33] n193 NOR2xp33_ASAP7_75t_R
XU1220 In_Weight[94] n1257 n192 NOR2xp33_ASAP7_75t_R
XU1221 weight_valid Weight[34] n195 NOR2xp33_ASAP7_75t_R
XU1222 In_Weight[93] n1257 n194 NOR2xp33_ASAP7_75t_R
XU1223 weight_valid Weight[35] n197 NOR2xp33_ASAP7_75t_R
XU1224 In_Weight[92] n1257 n196 NOR2xp33_ASAP7_75t_R
XU1225 weight_valid Weight[36] n199 NOR2xp33_ASAP7_75t_R
XU1226 In_Weight[91] n1258 n198 NOR2xp33_ASAP7_75t_R
XU1227 weight_valid Weight[37] n201 NOR2xp33_ASAP7_75t_R
XU1228 In_Weight[90] n1258 n200 NOR2xp33_ASAP7_75t_R
XU1229 weight_valid Weight[38] n203 NOR2xp33_ASAP7_75t_R
XU1230 In_Weight[89] n1258 n202 NOR2xp33_ASAP7_75t_R
XU1231 weight_valid Weight[39] n205 NOR2xp33_ASAP7_75t_R
XU1232 In_Weight[88] n1258 n204 NOR2xp33_ASAP7_75t_R
XU1233 weight_valid Weight[40] n207 NOR2xp33_ASAP7_75t_R
XU1234 In_Weight[87] n1258 n206 NOR2xp33_ASAP7_75t_R
XU1235 weight_valid Weight[41] n209 NOR2xp33_ASAP7_75t_R
XU1236 In_Weight[86] n1258 n208 NOR2xp33_ASAP7_75t_R
XU1237 weight_valid Weight[42] n211 NOR2xp33_ASAP7_75t_R
XU1238 In_Weight[85] n1258 n210 NOR2xp33_ASAP7_75t_R
XU1239 weight_valid Weight[43] n213 NOR2xp33_ASAP7_75t_R
XU1240 In_Weight[84] n1258 n212 NOR2xp33_ASAP7_75t_R
XU1241 weight_valid Weight[44] n215 NOR2xp33_ASAP7_75t_R
XU1242 In_Weight[83] n1258 n214 NOR2xp33_ASAP7_75t_R
XU1243 weight_valid Weight[45] n217 NOR2xp33_ASAP7_75t_R
XU1244 In_Weight[82] n1258 n216 NOR2xp33_ASAP7_75t_R
XU1245 weight_valid Weight[46] n219 NOR2xp33_ASAP7_75t_R
XU1246 In_Weight[81] n1258 n218 NOR2xp33_ASAP7_75t_R
XU1247 weight_valid Weight[47] n221 NOR2xp33_ASAP7_75t_R
XU1248 In_Weight[80] n1258 n220 NOR2xp33_ASAP7_75t_R
XU1249 weight_valid Weight[48] n223 NOR2xp33_ASAP7_75t_R
XU1250 In_Weight[79] n1259 n222 NOR2xp33_ASAP7_75t_R
XU1251 weight_valid Weight[49] n225 NOR2xp33_ASAP7_75t_R
XU1252 In_Weight[78] n1259 n224 NOR2xp33_ASAP7_75t_R
XU1253 weight_valid Weight[50] n227 NOR2xp33_ASAP7_75t_R
XU1254 In_Weight[77] n1259 n226 NOR2xp33_ASAP7_75t_R
XU1255 weight_valid Weight[51] n229 NOR2xp33_ASAP7_75t_R
XU1256 In_Weight[76] n1259 n228 NOR2xp33_ASAP7_75t_R
XU1257 weight_valid Weight[52] n231 NOR2xp33_ASAP7_75t_R
XU1258 In_Weight[75] n1259 n230 NOR2xp33_ASAP7_75t_R
XU1259 weight_valid Weight[53] n233 NOR2xp33_ASAP7_75t_R
XU1260 In_Weight[74] n1259 n232 NOR2xp33_ASAP7_75t_R
XU1261 weight_valid Weight[54] n235 NOR2xp33_ASAP7_75t_R
XU1262 In_Weight[73] n1259 n234 NOR2xp33_ASAP7_75t_R
XU1263 weight_valid Weight[55] n237 NOR2xp33_ASAP7_75t_R
XU1264 In_Weight[72] n1259 n236 NOR2xp33_ASAP7_75t_R
XU1265 weight_valid Weight[56] n239 NOR2xp33_ASAP7_75t_R
XU1266 In_Weight[71] n1259 n238 NOR2xp33_ASAP7_75t_R
XU1267 weight_valid Weight[57] n241 NOR2xp33_ASAP7_75t_R
XU1268 In_Weight[70] n1259 n240 NOR2xp33_ASAP7_75t_R
XU1269 weight_valid Weight[58] n243 NOR2xp33_ASAP7_75t_R
XU1270 In_Weight[69] n1259 n242 NOR2xp33_ASAP7_75t_R
XU1271 weight_valid Weight[59] n245 NOR2xp33_ASAP7_75t_R
XU1272 In_Weight[68] n1259 n244 NOR2xp33_ASAP7_75t_R
XU1273 weight_valid Weight[60] n247 NOR2xp33_ASAP7_75t_R
XU1274 In_Weight[67] n1260 n246 NOR2xp33_ASAP7_75t_R
XU1275 weight_valid Weight[61] n249 NOR2xp33_ASAP7_75t_R
XU1276 In_Weight[66] n1260 n248 NOR2xp33_ASAP7_75t_R
XU1277 weight_valid Weight[62] n251 NOR2xp33_ASAP7_75t_R
XU1278 In_Weight[65] n1260 n250 NOR2xp33_ASAP7_75t_R
XU1279 weight_valid Weight[63] n253 NOR2xp33_ASAP7_75t_R
XU1280 In_Weight[64] n1260 n252 NOR2xp33_ASAP7_75t_R
XU1281 weight_valid Weight[64] n255 NOR2xp33_ASAP7_75t_R
XU1282 In_Weight[63] n1260 n254 NOR2xp33_ASAP7_75t_R
XU1283 weight_valid Weight[65] n257 NOR2xp33_ASAP7_75t_R
XU1284 In_Weight[62] n1260 n256 NOR2xp33_ASAP7_75t_R
XU1285 weight_valid Weight[66] n259 NOR2xp33_ASAP7_75t_R
XU1286 In_Weight[61] n1260 n258 NOR2xp33_ASAP7_75t_R
XU1287 weight_valid Weight[67] n261 NOR2xp33_ASAP7_75t_R
XU1288 In_Weight[60] n1260 n260 NOR2xp33_ASAP7_75t_R
XU1289 weight_valid Weight[68] n263 NOR2xp33_ASAP7_75t_R
XU1290 In_Weight[59] n1260 n262 NOR2xp33_ASAP7_75t_R
XU1291 weight_valid Weight[69] n265 NOR2xp33_ASAP7_75t_R
XU1292 In_Weight[58] n1260 n264 NOR2xp33_ASAP7_75t_R
XU1293 weight_valid Weight[70] n267 NOR2xp33_ASAP7_75t_R
XU1294 In_Weight[57] n1260 n266 NOR2xp33_ASAP7_75t_R
XU1295 weight_valid Weight[71] n269 NOR2xp33_ASAP7_75t_R
XU1296 In_Weight[56] n1260 n268 NOR2xp33_ASAP7_75t_R
XU1297 weight_valid Weight[72] n271 NOR2xp33_ASAP7_75t_R
XU1298 In_Weight[55] n1259 n270 NOR2xp33_ASAP7_75t_R
XU1299 weight_valid Weight[73] n273 NOR2xp33_ASAP7_75t_R
XU1300 In_Weight[54] n1260 n272 NOR2xp33_ASAP7_75t_R
XU1301 weight_valid Weight[74] n275 NOR2xp33_ASAP7_75t_R
XU1302 In_Weight[53] n1255 n274 NOR2xp33_ASAP7_75t_R
XU1303 weight_valid Weight[75] n277 NOR2xp33_ASAP7_75t_R
XU1304 In_Weight[52] n1256 n276 NOR2xp33_ASAP7_75t_R
XU1305 weight_valid Weight[76] n279 NOR2xp33_ASAP7_75t_R
XU1306 In_Weight[51] n1257 n278 NOR2xp33_ASAP7_75t_R
XU1307 weight_valid Weight[77] n281 NOR2xp33_ASAP7_75t_R
XU1308 In_Weight[50] n1258 n280 NOR2xp33_ASAP7_75t_R
XU1309 weight_valid Weight[78] n283 NOR2xp33_ASAP7_75t_R
XU1310 In_Weight[49] n1259 n282 NOR2xp33_ASAP7_75t_R
XU1311 weight_valid Weight[79] n285 NOR2xp33_ASAP7_75t_R
XU1312 In_Weight[48] n1260 n284 NOR2xp33_ASAP7_75t_R
XU1313 weight_valid Weight[80] n287 NOR2xp33_ASAP7_75t_R
XU1314 In_Weight[47] n1255 n286 NOR2xp33_ASAP7_75t_R
XU1315 weight_valid Weight[81] n289 NOR2xp33_ASAP7_75t_R
XU1316 In_Weight[46] n1256 n288 NOR2xp33_ASAP7_75t_R
XU1317 weight_valid Weight[82] n291 NOR2xp33_ASAP7_75t_R
XU1318 In_Weight[45] n1257 n290 NOR2xp33_ASAP7_75t_R
XU1319 weight_valid Weight[83] n293 NOR2xp33_ASAP7_75t_R
XU1320 In_Weight[44] n1258 n292 NOR2xp33_ASAP7_75t_R
XU1321 weight_valid Weight[84] n295 NOR2xp33_ASAP7_75t_R
XU1322 In_Weight[43] n1258 n294 NOR2xp33_ASAP7_75t_R
XU1323 weight_valid Weight[85] n297 NOR2xp33_ASAP7_75t_R
XU1324 In_Weight[42] n1259 n296 NOR2xp33_ASAP7_75t_R
XU1325 weight_valid Weight[86] n299 NOR2xp33_ASAP7_75t_R
XU1326 In_Weight[41] n1256 n298 NOR2xp33_ASAP7_75t_R
XU1327 weight_valid Weight[87] n301 NOR2xp33_ASAP7_75t_R
XU1328 In_Weight[40] n1259 n300 NOR2xp33_ASAP7_75t_R
XU1329 weight_valid Weight[88] n303 NOR2xp33_ASAP7_75t_R
XU1330 In_Weight[39] n1260 n302 NOR2xp33_ASAP7_75t_R
XU1331 weight_valid Weight[89] n305 NOR2xp33_ASAP7_75t_R
XU1332 In_Weight[38] n1260 n304 NOR2xp33_ASAP7_75t_R
XU1333 weight_valid Weight[90] n307 NOR2xp33_ASAP7_75t_R
XU1334 In_Weight[37] n1257 n306 NOR2xp33_ASAP7_75t_R
XU1335 weight_valid Weight[91] n309 NOR2xp33_ASAP7_75t_R
XU1336 In_Weight[36] n1259 n308 NOR2xp33_ASAP7_75t_R
XU1337 weight_valid Weight[92] n311 NOR2xp33_ASAP7_75t_R
XU1338 In_Weight[35] n1255 n310 NOR2xp33_ASAP7_75t_R
XU1339 weight_valid Weight[93] n313 NOR2xp33_ASAP7_75t_R
XU1340 In_Weight[34] n1260 n312 NOR2xp33_ASAP7_75t_R
XU1341 weight_valid Weight[94] n315 NOR2xp33_ASAP7_75t_R
XU1342 In_Weight[33] n1258 n314 NOR2xp33_ASAP7_75t_R
XU1343 weight_valid Weight[95] n317 NOR2xp33_ASAP7_75t_R
XU1344 In_Weight[32] n1256 n316 NOR2xp33_ASAP7_75t_R
XU1345 weight_valid Weight[96] n319 NOR2xp33_ASAP7_75t_R
XU1346 In_Weight[31] n1258 n318 NOR2xp33_ASAP7_75t_R
XU1347 weight_valid Weight[97] n321 NOR2xp33_ASAP7_75t_R
XU1348 In_Weight[30] n1260 n320 NOR2xp33_ASAP7_75t_R
XU1349 weight_valid Weight[98] n323 NOR2xp33_ASAP7_75t_R
XU1350 In_Weight[29] n1257 n322 NOR2xp33_ASAP7_75t_R
XU1351 weight_valid Weight[99] n325 NOR2xp33_ASAP7_75t_R
XU1352 In_Weight[28] n1259 n324 NOR2xp33_ASAP7_75t_R
XU1353 weight_valid Weight[100] n327 NOR2xp33_ASAP7_75t_R
XU1354 In_Weight[27] n1260 n326 NOR2xp33_ASAP7_75t_R
XU1355 weight_valid Weight[101] n329 NOR2xp33_ASAP7_75t_R
XU1356 In_Weight[26] n1257 n328 NOR2xp33_ASAP7_75t_R
XU1357 weight_valid Weight[102] n331 NOR2xp33_ASAP7_75t_R
XU1358 In_Weight[25] n1258 n330 NOR2xp33_ASAP7_75t_R
XU1359 weight_valid Weight[103] n333 NOR2xp33_ASAP7_75t_R
XU1360 In_Weight[24] n1258 n332 NOR2xp33_ASAP7_75t_R
XU1361 weight_valid Weight[104] n335 NOR2xp33_ASAP7_75t_R
XU1362 In_Weight[23] n1255 n334 NOR2xp33_ASAP7_75t_R
XU1363 weight_valid Weight[105] n337 NOR2xp33_ASAP7_75t_R
XU1364 In_Weight[22] n1255 n336 NOR2xp33_ASAP7_75t_R
XU1365 weight_valid Weight[106] n339 NOR2xp33_ASAP7_75t_R
XU1366 In_Weight[21] n1259 n338 NOR2xp33_ASAP7_75t_R
XU1367 weight_valid Weight[107] n341 NOR2xp33_ASAP7_75t_R
XU1368 In_Weight[20] n1256 n340 NOR2xp33_ASAP7_75t_R
XU1369 weight_valid Weight[108] n343 NOR2xp33_ASAP7_75t_R
XU1370 In_Weight[19] n1259 n342 NOR2xp33_ASAP7_75t_R
XU1371 weight_valid Weight[109] n345 NOR2xp33_ASAP7_75t_R
XU1372 In_Weight[18] n1256 n344 NOR2xp33_ASAP7_75t_R
XU1373 weight_valid Weight[110] n347 NOR2xp33_ASAP7_75t_R
XU1374 In_Weight[17] n1255 n346 NOR2xp33_ASAP7_75t_R
XU1375 weight_valid Weight[111] n349 NOR2xp33_ASAP7_75t_R
XU1376 In_Weight[16] n1260 n348 NOR2xp33_ASAP7_75t_R
XU1377 weight_valid Weight[112] n351 NOR2xp33_ASAP7_75t_R
XU1378 In_Weight[15] n1257 n350 NOR2xp33_ASAP7_75t_R
XU1379 weight_valid Weight[113] n353 NOR2xp33_ASAP7_75t_R
XU1380 In_Weight[14] n1257 n352 NOR2xp33_ASAP7_75t_R
XU1381 weight_valid Weight[114] n355 NOR2xp33_ASAP7_75t_R
XU1382 In_Weight[13] n1256 n354 NOR2xp33_ASAP7_75t_R
XU1383 weight_valid Weight[115] n357 NOR2xp33_ASAP7_75t_R
XU1384 In_Weight[12] n1256 n356 NOR2xp33_ASAP7_75t_R
XU1385 weight_valid Weight[116] n359 NOR2xp33_ASAP7_75t_R
XU1386 In_Weight[11] n1257 n358 NOR2xp33_ASAP7_75t_R
XU1387 weight_valid Weight[117] n361 NOR2xp33_ASAP7_75t_R
XU1388 In_Weight[10] n1258 n360 NOR2xp33_ASAP7_75t_R
XU1389 weight_valid Weight[118] n363 NOR2xp33_ASAP7_75t_R
XU1390 In_Weight[9] n1255 n362 NOR2xp33_ASAP7_75t_R
XU1391 weight_valid Weight[119] n365 NOR2xp33_ASAP7_75t_R
XU1392 In_Weight[8] n1255 n364 NOR2xp33_ASAP7_75t_R
XU1393 in_valid n1261 INVx1_ASAP7_75t_R
XU1394 in_valid n1262 INVx1_ASAP7_75t_R
XU1395 in_valid n1263 INVx1_ASAP7_75t_R
XU1396 in_valid n1264 INVx1_ASAP7_75t_R
XU1397 in_valid n1265 INVx1_ASAP7_75t_R
XU1398 in_valid n1266 INVx1_ASAP7_75t_R
XU1399 in_valid IFM[0] n382 NOR2xp33_ASAP7_75t_R
XU1400 In_IFM[127] n1261 n383 NOR2xp33_ASAP7_75t_R
XU1401 in_valid IFM[1] n384 NOR2xp33_ASAP7_75t_R
XU1402 In_IFM[126] n1261 n385 NOR2xp33_ASAP7_75t_R
XU1403 in_valid IFM[2] n386 NOR2xp33_ASAP7_75t_R
XU1404 In_IFM[125] n1261 n387 NOR2xp33_ASAP7_75t_R
XU1405 in_valid IFM[3] n388 NOR2xp33_ASAP7_75t_R
XU1406 In_IFM[124] n1261 n389 NOR2xp33_ASAP7_75t_R
XU1407 in_valid IFM[4] n390 NOR2xp33_ASAP7_75t_R
XU1408 In_IFM[123] n1261 n391 NOR2xp33_ASAP7_75t_R
XU1409 in_valid IFM[5] n392 NOR2xp33_ASAP7_75t_R
XU1410 In_IFM[122] n1261 n393 NOR2xp33_ASAP7_75t_R
XU1411 in_valid IFM[6] n394 NOR2xp33_ASAP7_75t_R
XU1412 In_IFM[121] n1261 n395 NOR2xp33_ASAP7_75t_R
XU1413 in_valid IFM[7] n396 NOR2xp33_ASAP7_75t_R
XU1414 In_IFM[120] n1261 n397 NOR2xp33_ASAP7_75t_R
XU1415 in_valid IFM[8] n398 NOR2xp33_ASAP7_75t_R
XU1416 In_IFM[119] n1261 n399 NOR2xp33_ASAP7_75t_R
XU1417 in_valid IFM[9] n400 NOR2xp33_ASAP7_75t_R
XU1418 In_IFM[118] n1261 n401 NOR2xp33_ASAP7_75t_R
XU1419 in_valid IFM[10] n402 NOR2xp33_ASAP7_75t_R
XU1420 In_IFM[117] n1261 n403 NOR2xp33_ASAP7_75t_R
XU1421 in_valid IFM[11] n404 NOR2xp33_ASAP7_75t_R
XU1422 In_IFM[116] n1261 n405 NOR2xp33_ASAP7_75t_R
XU1423 in_valid IFM[12] n406 NOR2xp33_ASAP7_75t_R
XU1424 In_IFM[115] n1262 n407 NOR2xp33_ASAP7_75t_R
XU1425 in_valid IFM[13] n408 NOR2xp33_ASAP7_75t_R
XU1426 In_IFM[114] n1262 n409 NOR2xp33_ASAP7_75t_R
XU1427 in_valid IFM[14] n410 NOR2xp33_ASAP7_75t_R
XU1428 In_IFM[113] n1262 n411 NOR2xp33_ASAP7_75t_R
XU1429 in_valid IFM[15] n412 NOR2xp33_ASAP7_75t_R
XU1430 In_IFM[112] n1262 n413 NOR2xp33_ASAP7_75t_R
XU1431 in_valid IFM[16] n414 NOR2xp33_ASAP7_75t_R
XU1432 In_IFM[111] n1262 n415 NOR2xp33_ASAP7_75t_R
XU1433 in_valid IFM[17] n416 NOR2xp33_ASAP7_75t_R
XU1434 In_IFM[110] n1262 n417 NOR2xp33_ASAP7_75t_R
XU1435 in_valid IFM[18] n418 NOR2xp33_ASAP7_75t_R
XU1436 In_IFM[109] n1262 n419 NOR2xp33_ASAP7_75t_R
XU1437 in_valid IFM[19] n420 NOR2xp33_ASAP7_75t_R
XU1438 In_IFM[108] n1262 n421 NOR2xp33_ASAP7_75t_R
XU1439 in_valid IFM[20] n422 NOR2xp33_ASAP7_75t_R
XU1440 In_IFM[107] n1262 n423 NOR2xp33_ASAP7_75t_R
XU1441 in_valid IFM[21] n424 NOR2xp33_ASAP7_75t_R
XU1442 In_IFM[106] n1262 n425 NOR2xp33_ASAP7_75t_R
XU1443 in_valid IFM[22] n426 NOR2xp33_ASAP7_75t_R
XU1444 In_IFM[105] n1262 n427 NOR2xp33_ASAP7_75t_R
XU1445 in_valid IFM[23] n428 NOR2xp33_ASAP7_75t_R
XU1446 In_IFM[104] n1262 n429 NOR2xp33_ASAP7_75t_R
XU1447 in_valid IFM[24] n430 NOR2xp33_ASAP7_75t_R
XU1448 In_IFM[103] n1263 n431 NOR2xp33_ASAP7_75t_R
XU1449 in_valid IFM[25] n432 NOR2xp33_ASAP7_75t_R
XU1450 In_IFM[102] n1263 n433 NOR2xp33_ASAP7_75t_R
XU1451 in_valid IFM[26] n434 NOR2xp33_ASAP7_75t_R
XU1452 In_IFM[101] n1263 n435 NOR2xp33_ASAP7_75t_R
XU1453 in_valid IFM[27] n436 NOR2xp33_ASAP7_75t_R
XU1454 In_IFM[100] n1263 n437 NOR2xp33_ASAP7_75t_R
XU1455 in_valid IFM[28] n438 NOR2xp33_ASAP7_75t_R
XU1456 In_IFM[99] n1263 n439 NOR2xp33_ASAP7_75t_R
XU1457 in_valid IFM[29] n440 NOR2xp33_ASAP7_75t_R
XU1458 In_IFM[98] n1263 n441 NOR2xp33_ASAP7_75t_R
XU1459 in_valid IFM[30] n442 NOR2xp33_ASAP7_75t_R
XU1460 In_IFM[97] n1263 n443 NOR2xp33_ASAP7_75t_R
XU1461 in_valid IFM[31] n444 NOR2xp33_ASAP7_75t_R
XU1462 In_IFM[96] n1263 n445 NOR2xp33_ASAP7_75t_R
XU1463 in_valid IFM[32] n446 NOR2xp33_ASAP7_75t_R
XU1464 In_IFM[95] n1263 n447 NOR2xp33_ASAP7_75t_R
XU1465 in_valid IFM[33] n448 NOR2xp33_ASAP7_75t_R
XU1466 In_IFM[94] n1263 n449 NOR2xp33_ASAP7_75t_R
XU1467 in_valid IFM[34] n450 NOR2xp33_ASAP7_75t_R
XU1468 In_IFM[93] n1263 n451 NOR2xp33_ASAP7_75t_R
XU1469 in_valid IFM[35] n452 NOR2xp33_ASAP7_75t_R
XU1470 In_IFM[92] n1263 n453 NOR2xp33_ASAP7_75t_R
XU1471 in_valid IFM[36] n454 NOR2xp33_ASAP7_75t_R
XU1472 In_IFM[91] n1264 n455 NOR2xp33_ASAP7_75t_R
XU1473 in_valid IFM[37] n456 NOR2xp33_ASAP7_75t_R
XU1474 In_IFM[90] n1264 n457 NOR2xp33_ASAP7_75t_R
XU1475 in_valid IFM[38] n458 NOR2xp33_ASAP7_75t_R
XU1476 In_IFM[89] n1264 n459 NOR2xp33_ASAP7_75t_R
XU1477 in_valid IFM[39] n460 NOR2xp33_ASAP7_75t_R
XU1478 In_IFM[88] n1264 n461 NOR2xp33_ASAP7_75t_R
XU1479 in_valid IFM[40] n462 NOR2xp33_ASAP7_75t_R
XU1480 In_IFM[87] n1264 n463 NOR2xp33_ASAP7_75t_R
XU1481 in_valid IFM[41] n464 NOR2xp33_ASAP7_75t_R
XU1482 In_IFM[86] n1264 n465 NOR2xp33_ASAP7_75t_R
XU1483 in_valid IFM[42] n466 NOR2xp33_ASAP7_75t_R
XU1484 In_IFM[85] n1264 n467 NOR2xp33_ASAP7_75t_R
XU1485 in_valid IFM[43] n468 NOR2xp33_ASAP7_75t_R
XU1486 In_IFM[84] n1264 n469 NOR2xp33_ASAP7_75t_R
XU1487 in_valid IFM[44] n470 NOR2xp33_ASAP7_75t_R
XU1488 In_IFM[83] n1264 n471 NOR2xp33_ASAP7_75t_R
XU1489 in_valid IFM[45] n472 NOR2xp33_ASAP7_75t_R
XU1490 In_IFM[82] n1264 n473 NOR2xp33_ASAP7_75t_R
XU1491 in_valid IFM[46] n474 NOR2xp33_ASAP7_75t_R
XU1492 In_IFM[81] n1264 n475 NOR2xp33_ASAP7_75t_R
XU1493 in_valid IFM[47] n476 NOR2xp33_ASAP7_75t_R
XU1494 In_IFM[80] n1264 n477 NOR2xp33_ASAP7_75t_R
XU1495 in_valid IFM[48] n478 NOR2xp33_ASAP7_75t_R
XU1496 In_IFM[79] n1265 n479 NOR2xp33_ASAP7_75t_R
XU1497 in_valid IFM[49] n480 NOR2xp33_ASAP7_75t_R
XU1498 In_IFM[78] n1265 n481 NOR2xp33_ASAP7_75t_R
XU1499 in_valid IFM[50] n482 NOR2xp33_ASAP7_75t_R
XU1500 In_IFM[77] n1265 n483 NOR2xp33_ASAP7_75t_R
XU1501 in_valid IFM[51] n484 NOR2xp33_ASAP7_75t_R
XU1502 In_IFM[76] n1265 n485 NOR2xp33_ASAP7_75t_R
XU1503 in_valid IFM[52] n486 NOR2xp33_ASAP7_75t_R
XU1504 In_IFM[75] n1265 n487 NOR2xp33_ASAP7_75t_R
XU1505 in_valid IFM[53] n488 NOR2xp33_ASAP7_75t_R
XU1506 In_IFM[74] n1265 n489 NOR2xp33_ASAP7_75t_R
XU1507 in_valid IFM[54] n490 NOR2xp33_ASAP7_75t_R
XU1508 In_IFM[73] n1265 n491 NOR2xp33_ASAP7_75t_R
XU1509 in_valid IFM[55] n492 NOR2xp33_ASAP7_75t_R
XU1510 In_IFM[72] n1265 n493 NOR2xp33_ASAP7_75t_R
XU1511 in_valid IFM[56] n494 NOR2xp33_ASAP7_75t_R
XU1512 In_IFM[71] n1265 n495 NOR2xp33_ASAP7_75t_R
XU1513 in_valid IFM[57] n496 NOR2xp33_ASAP7_75t_R
XU1514 In_IFM[70] n1265 n497 NOR2xp33_ASAP7_75t_R
XU1515 in_valid IFM[58] n498 NOR2xp33_ASAP7_75t_R
XU1516 In_IFM[69] n1265 n499 NOR2xp33_ASAP7_75t_R
XU1517 in_valid IFM[59] n500 NOR2xp33_ASAP7_75t_R
XU1518 In_IFM[68] n1265 n501 NOR2xp33_ASAP7_75t_R
XU1519 in_valid IFM[60] n502 NOR2xp33_ASAP7_75t_R
XU1520 In_IFM[67] n1266 n503 NOR2xp33_ASAP7_75t_R
XU1521 in_valid IFM[61] n504 NOR2xp33_ASAP7_75t_R
XU1522 In_IFM[66] n1266 n505 NOR2xp33_ASAP7_75t_R
XU1523 in_valid IFM[62] n506 NOR2xp33_ASAP7_75t_R
XU1524 In_IFM[65] n1266 n507 NOR2xp33_ASAP7_75t_R
XU1525 in_valid IFM[63] n508 NOR2xp33_ASAP7_75t_R
XU1526 In_IFM[64] n1266 n509 NOR2xp33_ASAP7_75t_R
XU1527 in_valid IFM[64] n510 NOR2xp33_ASAP7_75t_R
XU1528 In_IFM[63] n1266 n511 NOR2xp33_ASAP7_75t_R
XU1529 in_valid IFM[65] n512 NOR2xp33_ASAP7_75t_R
XU1530 In_IFM[62] n1266 n513 NOR2xp33_ASAP7_75t_R
XU1531 in_valid IFM[66] n514 NOR2xp33_ASAP7_75t_R
XU1532 In_IFM[61] n1266 n515 NOR2xp33_ASAP7_75t_R
XU1533 in_valid IFM[67] n516 NOR2xp33_ASAP7_75t_R
XU1534 In_IFM[60] n1266 n517 NOR2xp33_ASAP7_75t_R
XU1535 in_valid IFM[68] n518 NOR2xp33_ASAP7_75t_R
XU1536 In_IFM[59] n1266 n519 NOR2xp33_ASAP7_75t_R
XU1537 in_valid IFM[69] n520 NOR2xp33_ASAP7_75t_R
XU1538 In_IFM[58] n1266 n521 NOR2xp33_ASAP7_75t_R
XU1539 in_valid IFM[70] n522 NOR2xp33_ASAP7_75t_R
XU1540 In_IFM[57] n1266 n523 NOR2xp33_ASAP7_75t_R
XU1541 in_valid IFM[71] n524 NOR2xp33_ASAP7_75t_R
XU1542 In_IFM[56] n1266 n525 NOR2xp33_ASAP7_75t_R
XU1543 in_valid IFM[72] n526 NOR2xp33_ASAP7_75t_R
XU1544 In_IFM[55] n1263 n527 NOR2xp33_ASAP7_75t_R
XU1545 in_valid IFM[73] n528 NOR2xp33_ASAP7_75t_R
XU1546 In_IFM[54] n1264 n529 NOR2xp33_ASAP7_75t_R
XU1547 in_valid IFM[74] n530 NOR2xp33_ASAP7_75t_R
XU1548 In_IFM[53] n1261 n531 NOR2xp33_ASAP7_75t_R
XU1549 in_valid IFM[75] n532 NOR2xp33_ASAP7_75t_R
XU1550 In_IFM[52] n1265 n533 NOR2xp33_ASAP7_75t_R
XU1551 in_valid IFM[76] n534 NOR2xp33_ASAP7_75t_R
XU1552 In_IFM[51] n1266 n535 NOR2xp33_ASAP7_75t_R
XU1553 in_valid IFM[77] n536 NOR2xp33_ASAP7_75t_R
XU1554 In_IFM[50] n1262 n537 NOR2xp33_ASAP7_75t_R
XU1555 in_valid IFM[78] n538 NOR2xp33_ASAP7_75t_R
XU1556 In_IFM[49] n1263 n539 NOR2xp33_ASAP7_75t_R
XU1557 in_valid IFM[79] n540 NOR2xp33_ASAP7_75t_R
XU1558 In_IFM[48] n1264 n541 NOR2xp33_ASAP7_75t_R
XU1559 in_valid IFM[80] n542 NOR2xp33_ASAP7_75t_R
XU1560 In_IFM[47] n1261 n543 NOR2xp33_ASAP7_75t_R
XU1561 in_valid IFM[81] n544 NOR2xp33_ASAP7_75t_R
XU1562 In_IFM[46] n1265 n545 NOR2xp33_ASAP7_75t_R
XU1563 in_valid IFM[82] n546 NOR2xp33_ASAP7_75t_R
XU1564 In_IFM[45] n1266 n547 NOR2xp33_ASAP7_75t_R
XU1565 in_valid IFM[83] n548 NOR2xp33_ASAP7_75t_R
XU1566 In_IFM[44] n1262 n549 NOR2xp33_ASAP7_75t_R
XU1567 in_valid IFM[84] n550 NOR2xp33_ASAP7_75t_R
XU1568 In_IFM[43] n1265 n551 NOR2xp33_ASAP7_75t_R
XU1569 in_valid IFM[85] n552 NOR2xp33_ASAP7_75t_R
XU1570 In_IFM[42] n1261 n553 NOR2xp33_ASAP7_75t_R
XU1571 in_valid IFM[86] n554 NOR2xp33_ASAP7_75t_R
XU1572 In_IFM[41] n1262 n555 NOR2xp33_ASAP7_75t_R
XU1573 in_valid IFM[87] n556 NOR2xp33_ASAP7_75t_R
XU1574 In_IFM[40] n1263 n557 NOR2xp33_ASAP7_75t_R
XU1575 in_valid IFM[88] n558 NOR2xp33_ASAP7_75t_R
XU1576 In_IFM[39] n1264 n559 NOR2xp33_ASAP7_75t_R
XU1577 in_valid IFM[89] n560 NOR2xp33_ASAP7_75t_R
XU1578 In_IFM[38] n1265 n561 NOR2xp33_ASAP7_75t_R
XU1579 in_valid IFM[90] n562 NOR2xp33_ASAP7_75t_R
XU1580 In_IFM[37] n1266 n563 NOR2xp33_ASAP7_75t_R
XU1581 in_valid IFM[91] n564 NOR2xp33_ASAP7_75t_R
XU1582 In_IFM[36] n1266 n565 NOR2xp33_ASAP7_75t_R
XU1583 in_valid IFM[92] n566 NOR2xp33_ASAP7_75t_R
XU1584 In_IFM[35] n1261 n567 NOR2xp33_ASAP7_75t_R
XU1585 in_valid IFM[93] n568 NOR2xp33_ASAP7_75t_R
XU1586 In_IFM[34] n1262 n569 NOR2xp33_ASAP7_75t_R
XU1587 in_valid IFM[94] n570 NOR2xp33_ASAP7_75t_R
XU1588 In_IFM[33] n1263 n571 NOR2xp33_ASAP7_75t_R
XU1589 in_valid IFM[95] n572 NOR2xp33_ASAP7_75t_R
XU1590 In_IFM[32] n1264 n573 NOR2xp33_ASAP7_75t_R
XU1591 in_valid IFM[96] n574 NOR2xp33_ASAP7_75t_R
XU1592 In_IFM[31] n1261 n575 NOR2xp33_ASAP7_75t_R
XU1593 in_valid IFM[97] n576 NOR2xp33_ASAP7_75t_R
XU1594 In_IFM[30] n1262 n577 NOR2xp33_ASAP7_75t_R
XU1595 in_valid IFM[98] n578 NOR2xp33_ASAP7_75t_R
XU1596 In_IFM[29] n1261 n579 NOR2xp33_ASAP7_75t_R
XU1597 in_valid IFM[99] n580 NOR2xp33_ASAP7_75t_R
XU1598 In_IFM[28] n1266 n581 NOR2xp33_ASAP7_75t_R
XU1599 in_valid IFM[100] n582 NOR2xp33_ASAP7_75t_R
XU1600 In_IFM[27] n1265 n583 NOR2xp33_ASAP7_75t_R
XU1601 in_valid IFM[101] n584 NOR2xp33_ASAP7_75t_R
XU1602 In_IFM[26] n1263 n585 NOR2xp33_ASAP7_75t_R
XU1603 in_valid IFM[102] n586 NOR2xp33_ASAP7_75t_R
XU1604 In_IFM[25] n1265 n587 NOR2xp33_ASAP7_75t_R
XU1605 in_valid IFM[103] n588 NOR2xp33_ASAP7_75t_R
XU1606 In_IFM[24] n1262 n589 NOR2xp33_ASAP7_75t_R
XU1607 in_valid IFM[104] n590 NOR2xp33_ASAP7_75t_R
XU1608 In_IFM[23] n1263 n591 NOR2xp33_ASAP7_75t_R
XU1609 in_valid IFM[105] n592 NOR2xp33_ASAP7_75t_R
XU1610 In_IFM[22] n1264 n593 NOR2xp33_ASAP7_75t_R
XU1611 in_valid IFM[106] n594 NOR2xp33_ASAP7_75t_R
XU1612 In_IFM[21] n1261 n595 NOR2xp33_ASAP7_75t_R
XU1613 in_valid IFM[107] n596 NOR2xp33_ASAP7_75t_R
XU1614 In_IFM[20] n1266 n597 NOR2xp33_ASAP7_75t_R
XU1615 in_valid IFM[108] n598 NOR2xp33_ASAP7_75t_R
XU1616 In_IFM[19] n1262 n599 NOR2xp33_ASAP7_75t_R
XU1617 in_valid IFM[109] n600 NOR2xp33_ASAP7_75t_R
XU1618 In_IFM[18] n1263 n601 NOR2xp33_ASAP7_75t_R
XU1619 in_valid IFM[110] n602 NOR2xp33_ASAP7_75t_R
XU1620 In_IFM[17] n1264 n603 NOR2xp33_ASAP7_75t_R
XU1621 in_valid IFM[111] n604 NOR2xp33_ASAP7_75t_R
XU1622 In_IFM[16] n1265 n605 NOR2xp33_ASAP7_75t_R
XU1623 in_valid IFM[112] n606 NOR2xp33_ASAP7_75t_R
XU1624 In_IFM[15] n1266 n607 NOR2xp33_ASAP7_75t_R
XU1625 in_valid IFM[113] n608 NOR2xp33_ASAP7_75t_R
XU1626 In_IFM[14] n1266 n609 NOR2xp33_ASAP7_75t_R
XU1627 in_valid IFM[114] n610 NOR2xp33_ASAP7_75t_R
XU1628 In_IFM[13] n1264 n611 NOR2xp33_ASAP7_75t_R
XU1629 in_valid IFM[115] n612 NOR2xp33_ASAP7_75t_R
XU1630 In_IFM[12] n1266 n613 NOR2xp33_ASAP7_75t_R
XU1631 in_valid IFM[116] n614 NOR2xp33_ASAP7_75t_R
XU1632 In_IFM[11] n1261 n615 NOR2xp33_ASAP7_75t_R
XU1633 in_valid IFM[117] n616 NOR2xp33_ASAP7_75t_R
XU1634 In_IFM[10] n1262 n617 NOR2xp33_ASAP7_75t_R
XU1635 in_valid IFM[118] n618 NOR2xp33_ASAP7_75t_R
XU1636 In_IFM[9] n1263 n619 NOR2xp33_ASAP7_75t_R
XU1637 in_valid IFM[119] n620 NOR2xp33_ASAP7_75t_R
XU1638 In_IFM[8] n1264 n621 NOR2xp33_ASAP7_75t_R
XU1639 weight_valid Weight[120] n367 NOR2xp33_ASAP7_75t_R
XU1640 In_Weight[7] n1259 n366 NOR2xp33_ASAP7_75t_R
XU1641 weight_valid Weight[121] n369 NOR2xp33_ASAP7_75t_R
XU1642 In_Weight[6] n1257 n368 NOR2xp33_ASAP7_75t_R
XU1643 weight_valid Weight[122] n371 NOR2xp33_ASAP7_75t_R
XU1644 In_Weight[5] n1255 n370 NOR2xp33_ASAP7_75t_R
XU1645 weight_valid Weight[123] n373 NOR2xp33_ASAP7_75t_R
XU1646 In_Weight[4] n1260 n372 NOR2xp33_ASAP7_75t_R
XU1647 weight_valid Weight[124] n375 NOR2xp33_ASAP7_75t_R
XU1648 In_Weight[3] n1258 n374 NOR2xp33_ASAP7_75t_R
XU1649 weight_valid Weight[125] n377 NOR2xp33_ASAP7_75t_R
XU1650 In_Weight[2] n1258 n376 NOR2xp33_ASAP7_75t_R
XU1651 weight_valid Weight[126] n379 NOR2xp33_ASAP7_75t_R
XU1652 In_Weight[1] n1256 n378 NOR2xp33_ASAP7_75t_R
XU1653 weight_valid Weight[127] n381 NOR2xp33_ASAP7_75t_R
XU1654 In_Weight[0] n1257 n380 NOR2xp33_ASAP7_75t_R
XU1655 in_valid IFM[120] n622 NOR2xp33_ASAP7_75t_R
XU1656 In_IFM[7] n1262 n623 NOR2xp33_ASAP7_75t_R
XU1657 in_valid IFM[121] n624 NOR2xp33_ASAP7_75t_R
XU1658 In_IFM[6] n1263 n625 NOR2xp33_ASAP7_75t_R
XU1659 in_valid IFM[122] n626 NOR2xp33_ASAP7_75t_R
XU1660 In_IFM[5] n1264 n627 NOR2xp33_ASAP7_75t_R
XU1661 in_valid IFM[123] n628 NOR2xp33_ASAP7_75t_R
XU1662 In_IFM[4] n1265 n629 NOR2xp33_ASAP7_75t_R
XU1663 in_valid IFM[124] n630 NOR2xp33_ASAP7_75t_R
XU1664 In_IFM[3] n1266 n631 NOR2xp33_ASAP7_75t_R
XU1665 in_valid IFM[125] n632 NOR2xp33_ASAP7_75t_R
XU1666 In_IFM[2] n1262 n633 NOR2xp33_ASAP7_75t_R
XU1667 in_valid IFM[126] n634 NOR2xp33_ASAP7_75t_R
XU1668 In_IFM[1] n1265 n635 NOR2xp33_ASAP7_75t_R
XU1669 in_valid IFM[127] n636 NOR2xp33_ASAP7_75t_R
XU1670 In_IFM[0] n1265 n637 NOR2xp33_ASAP7_75t_R
XU1671 clk21 n1269 HB1xp67_ASAP7_75t_R
XU1672 clk21 rst_n n1267 AND2x2_ASAP7_75t_R
XU1673 rst_n n1270 n1268 AND2x4_ASAP7_75t_R
XU1674 N1308 state_cs n668 NAND2xp5_ASAP7_75t_R
XU1675 clk21 n1270 INVx1_ASAP7_75t_R
XU1676 Out_OFM2[0] n1268 n1272 NAND2xp5_ASAP7_75t_R
XU1677 n1267 Out_OFM1[0] n1271 NAND2xp5_ASAP7_75t_R
XU1678 n1272 n1271 Out_OFM[0] NAND2xp5_ASAP7_75t_R
XU1679 N1309 state_cs n669 NAND2xp5_ASAP7_75t_R
XU1680 Out_OFM2[1] n1268 n1274 NAND2xp5_ASAP7_75t_R
XU1681 n1267 Out_OFM1[1] n1273 NAND2xp5_ASAP7_75t_R
XU1682 n1274 n1273 Out_OFM[1] NAND2xp5_ASAP7_75t_R
XU1683 N1310 state_cs n670 NAND2xp5_ASAP7_75t_R
XU1684 Out_OFM2[2] n1268 n1276 NAND2xp5_ASAP7_75t_R
XU1685 n1267 Out_OFM1[2] n1275 NAND2xp5_ASAP7_75t_R
XU1686 n1276 n1275 Out_OFM[2] NAND2xp5_ASAP7_75t_R
XU1687 N1311 state_cs n671 NAND2xp5_ASAP7_75t_R
XU1688 Out_OFM2[3] n1268 n1278 NAND2xp5_ASAP7_75t_R
XU1689 n1267 Out_OFM1[3] n1277 NAND2xp5_ASAP7_75t_R
XU1690 n1278 n1277 Out_OFM[3] NAND2xp5_ASAP7_75t_R
XU1691 N1312 state_cs n672 NAND2xp5_ASAP7_75t_R
XU1692 Out_OFM2[4] n1268 n1280 NAND2xp5_ASAP7_75t_R
XU1693 n1267 Out_OFM1[4] n1279 NAND2xp5_ASAP7_75t_R
XU1694 n1280 n1279 Out_OFM[4] NAND2xp5_ASAP7_75t_R
XU1695 N1313 state_cs n673 NAND2xp5_ASAP7_75t_R
XU1696 Out_OFM2[5] n1268 n1282 NAND2xp5_ASAP7_75t_R
XU1697 n1267 Out_OFM1[5] n1281 NAND2xp5_ASAP7_75t_R
XU1698 n1282 n1281 Out_OFM[5] NAND2xp5_ASAP7_75t_R
XU1699 N1314 state_cs n674 NAND2xp5_ASAP7_75t_R
XU1700 Out_OFM2[6] n1268 n1284 NAND2xp5_ASAP7_75t_R
XU1701 n1267 Out_OFM1[6] n1283 NAND2xp5_ASAP7_75t_R
XU1702 n1284 n1283 Out_OFM[6] NAND2xp5_ASAP7_75t_R
XU1703 N1315 state_cs n675 NAND2xp5_ASAP7_75t_R
XU1704 Out_OFM2[7] n1268 n1286 NAND2xp5_ASAP7_75t_R
XU1705 n1267 Out_OFM1[7] n1285 NAND2xp5_ASAP7_75t_R
XU1706 n1286 n1285 Out_OFM[7] NAND2xp5_ASAP7_75t_R
XU1707 N1316 state_cs n676 NAND2xp5_ASAP7_75t_R
XU1708 Out_OFM2[8] n1268 n1288 NAND2xp5_ASAP7_75t_R
XU1709 n1267 Out_OFM1[8] n1287 NAND2xp5_ASAP7_75t_R
XU1710 n1288 n1287 Out_OFM[8] NAND2xp5_ASAP7_75t_R
XU1711 N1317 state_cs n677 NAND2xp5_ASAP7_75t_R
XU1712 Out_OFM2[9] n1268 n1290 NAND2xp5_ASAP7_75t_R
XU1713 Out_OFM1[9] n1267 n1289 NAND2xp5_ASAP7_75t_R
XU1714 n1290 n1289 Out_OFM[9] NAND2xp5_ASAP7_75t_R
XU1715 N1318 state_cs n678 NAND2xp5_ASAP7_75t_R
XU1716 Out_OFM2[10] n1268 n1292 NAND2xp5_ASAP7_75t_R
XU1717 n1267 Out_OFM1[10] n1291 NAND2xp5_ASAP7_75t_R
XU1718 n1292 n1291 Out_OFM[10] NAND2xp5_ASAP7_75t_R
XU1719 N1319 state_cs n679 NAND2xp5_ASAP7_75t_R
XU1720 Out_OFM2[11] n1268 n1294 NAND2xp5_ASAP7_75t_R
XU1721 Out_OFM1[11] n1267 n1293 NAND2xp5_ASAP7_75t_R
XU1722 n1294 n1293 Out_OFM[11] NAND2xp5_ASAP7_75t_R
XU1723 N1320 state_cs n680 NAND2xp5_ASAP7_75t_R
XU1724 Out_OFM2[12] n1268 n1296 NAND2xp5_ASAP7_75t_R
XU1725 n1267 Out_OFM1[12] n1295 NAND2xp5_ASAP7_75t_R
XU1726 n1296 n1295 Out_OFM[12] NAND2xp5_ASAP7_75t_R
XU1727 n1297 N1141 INVx1_ASAP7_75t_R
XU1728 n1299 N1142 INVx1_ASAP7_75t_R
XU1729 n1301 N1143 INVx1_ASAP7_75t_R
XU1730 n1303 N1144 INVx1_ASAP7_75t_R
XU1731 n1305 N1145 INVx1_ASAP7_75t_R
XU1732 n1307 N1146 INVx1_ASAP7_75t_R
XU1733 n1309 N1147 INVx1_ASAP7_75t_R
XU1734 n1310 N1148 INVx1_ASAP7_75t_R
XU1735 n1298 n1311 INVx1_ASAP7_75t_R
XU1736 n1300 n1312 INVx1_ASAP7_75t_R
XU1737 n1302 n1313 INVx1_ASAP7_75t_R
XU1738 n1304 n1314 INVx1_ASAP7_75t_R
XU1739 n1306 n1315 INVx1_ASAP7_75t_R
XU1740 n1308 n1316 INVx1_ASAP7_75t_R
XU1741 n1317 N1288 INVx1_ASAP7_75t_R
XU1742 n1319 N1289 INVx1_ASAP7_75t_R
XU1743 n1321 N1290 INVx1_ASAP7_75t_R
XU1744 n1323 N1291 INVx1_ASAP7_75t_R
XU1745 n1325 N1292 INVx1_ASAP7_75t_R
XU1746 n1327 N1293 INVx1_ASAP7_75t_R
XU1747 n1329 N1294 INVx1_ASAP7_75t_R
XU1748 n1330 N1295 INVx1_ASAP7_75t_R
XU1749 n1318 n1331 INVx1_ASAP7_75t_R
XU1750 n1320 n1332 INVx1_ASAP7_75t_R
XU1751 n1322 n1333 INVx1_ASAP7_75t_R
XU1752 n1324 n1334 INVx1_ASAP7_75t_R
XU1753 n1326 n1335 INVx1_ASAP7_75t_R
XU1754 n1328 n1336 INVx1_ASAP7_75t_R
XU1755 n1337 N1078 INVx1_ASAP7_75t_R
XU1756 n1339 N1079 INVx1_ASAP7_75t_R
XU1757 n1341 N1080 INVx1_ASAP7_75t_R
XU1758 n1343 N1081 INVx1_ASAP7_75t_R
XU1759 n1345 N1082 INVx1_ASAP7_75t_R
XU1760 n1347 N1083 INVx1_ASAP7_75t_R
XU1761 n1349 N1084 INVx1_ASAP7_75t_R
XU1762 n1351 N1085 INVx1_ASAP7_75t_R
XU1763 n1352 N1086 INVx1_ASAP7_75t_R
XU1764 n1338 n1353 INVx1_ASAP7_75t_R
XU1765 n1340 n1354 INVx1_ASAP7_75t_R
XU1766 n1342 n1355 INVx1_ASAP7_75t_R
XU1767 n1344 n1356 INVx1_ASAP7_75t_R
XU1768 n1346 n1357 INVx1_ASAP7_75t_R
XU1769 n1348 n1358 INVx1_ASAP7_75t_R
XU1770 n1350 n1359 INVx1_ASAP7_75t_R
XU1771 n1360 N994 INVx1_ASAP7_75t_R
XU1772 n1362 N995 INVx1_ASAP7_75t_R
XU1773 n1364 N996 INVx1_ASAP7_75t_R
XU1774 n1366 N997 INVx1_ASAP7_75t_R
XU1775 n1368 N998 INVx1_ASAP7_75t_R
XU1776 n1370 N999 INVx1_ASAP7_75t_R
XU1777 n1372 N1000 INVx1_ASAP7_75t_R
XU1778 n1373 N1001 INVx1_ASAP7_75t_R
XU1779 n1361 n1374 INVx1_ASAP7_75t_R
XU1780 n1363 n1375 INVx1_ASAP7_75t_R
XU1781 n1365 n1376 INVx1_ASAP7_75t_R
XU1782 n1367 n1377 INVx1_ASAP7_75t_R
XU1783 n1369 n1378 INVx1_ASAP7_75t_R
XU1784 n1371 n1379 INVx1_ASAP7_75t_R
XU1785 n1380 N910 INVx1_ASAP7_75t_R
XU1786 n1382 N911 INVx1_ASAP7_75t_R
XU1787 n1384 N912 INVx1_ASAP7_75t_R
XU1788 n1386 N913 INVx1_ASAP7_75t_R
XU1789 n1388 N914 INVx1_ASAP7_75t_R
XU1790 n1390 N915 INVx1_ASAP7_75t_R
XU1791 n1392 N916 INVx1_ASAP7_75t_R
XU1792 n1393 N917 INVx1_ASAP7_75t_R
XU1793 n1381 n1394 INVx1_ASAP7_75t_R
XU1794 n1383 n1395 INVx1_ASAP7_75t_R
XU1795 n1385 n1396 INVx1_ASAP7_75t_R
XU1796 n1387 n1397 INVx1_ASAP7_75t_R
XU1797 n1389 n1398 INVx1_ASAP7_75t_R
XU1798 n1391 n1399 INVx1_ASAP7_75t_R
XU1799 n1400 add_5_root_r893_B_1_ INVx1_ASAP7_75t_R
XU1800 n1402 add_5_root_r893_B_2_ INVx1_ASAP7_75t_R
XU1801 n1404 add_5_root_r893_B_3_ INVx1_ASAP7_75t_R
XU1802 n1406 add_5_root_r893_B_4_ INVx1_ASAP7_75t_R
XU1803 n1408 add_5_root_r893_B_5_ INVx1_ASAP7_75t_R
XU1804 n1410 add_5_root_r893_B_6_ INVx1_ASAP7_75t_R
XU1805 n1412 add_5_root_r893_B_7_ INVx1_ASAP7_75t_R
XU1806 n1414 add_5_root_r893_B_8_ INVx1_ASAP7_75t_R
XU1807 n1415 add_5_root_r893_B_9_ INVx1_ASAP7_75t_R
XU1808 n1401 n1416 INVx1_ASAP7_75t_R
XU1809 n1403 n1417 INVx1_ASAP7_75t_R
XU1810 n1405 n1418 INVx1_ASAP7_75t_R
XU1811 n1407 n1419 INVx1_ASAP7_75t_R
XU1812 n1409 n1420 INVx1_ASAP7_75t_R
XU1813 n1411 n1421 INVx1_ASAP7_75t_R
XU1814 n1413 n1422 INVx1_ASAP7_75t_R
XU1815 n1440 add_5_root_r893_SUM_10_ INVx1_ASAP7_75t_R
XU1816 n1423 add_5_root_r893_SUM_1_ INVx1_ASAP7_75t_R
XU1817 n1425 add_5_root_r893_SUM_2_ INVx1_ASAP7_75t_R
XU1818 n1427 add_5_root_r893_SUM_3_ INVx1_ASAP7_75t_R
XU1819 n1429 add_5_root_r893_SUM_4_ INVx1_ASAP7_75t_R
XU1820 n1431 add_5_root_r893_SUM_5_ INVx1_ASAP7_75t_R
XU1821 n1433 add_5_root_r893_SUM_6_ INVx1_ASAP7_75t_R
XU1822 n1435 add_5_root_r893_SUM_7_ INVx1_ASAP7_75t_R
XU1823 n1437 add_5_root_r893_SUM_8_ INVx1_ASAP7_75t_R
XU1824 n1439 add_5_root_r893_SUM_9_ INVx1_ASAP7_75t_R
XU1825 n1424 n1441 INVx1_ASAP7_75t_R
XU1826 n1426 n1442 INVx1_ASAP7_75t_R
XU1827 n1428 n1443 INVx1_ASAP7_75t_R
XU1828 n1430 n1444 INVx1_ASAP7_75t_R
XU1829 n1432 n1445 INVx1_ASAP7_75t_R
XU1830 n1434 n1446 INVx1_ASAP7_75t_R
XU1831 n1436 n1447 INVx1_ASAP7_75t_R
XU1832 n1438 n1448 INVx1_ASAP7_75t_R
XU1833 n1449 N952 INVx1_ASAP7_75t_R
XU1834 n1451 N953 INVx1_ASAP7_75t_R
XU1835 n1453 N954 INVx1_ASAP7_75t_R
XU1836 n1455 N955 INVx1_ASAP7_75t_R
XU1837 n1457 N956 INVx1_ASAP7_75t_R
XU1838 n1459 N957 INVx1_ASAP7_75t_R
XU1839 n1461 N958 INVx1_ASAP7_75t_R
XU1840 n1462 N959 INVx1_ASAP7_75t_R
XU1841 n1450 n1463 INVx1_ASAP7_75t_R
XU1842 n1452 n1464 INVx1_ASAP7_75t_R
XU1843 n1454 n1465 INVx1_ASAP7_75t_R
XU1844 n1456 n1466 INVx1_ASAP7_75t_R
XU1845 n1458 n1467 INVx1_ASAP7_75t_R
XU1846 n1460 n1468 INVx1_ASAP7_75t_R
XU1847 n1469 N1162 INVx1_ASAP7_75t_R
XU1848 n1471 N1163 INVx1_ASAP7_75t_R
XU1849 n1473 N1164 INVx1_ASAP7_75t_R
XU1850 n1475 N1165 INVx1_ASAP7_75t_R
XU1851 n1477 N1166 INVx1_ASAP7_75t_R
XU1852 n1479 N1167 INVx1_ASAP7_75t_R
XU1853 n1481 N1168 INVx1_ASAP7_75t_R
XU1854 n1482 N1169 INVx1_ASAP7_75t_R
XU1855 n1470 n1483 INVx1_ASAP7_75t_R
XU1856 n1472 n1484 INVx1_ASAP7_75t_R
XU1857 n1474 n1485 INVx1_ASAP7_75t_R
XU1858 n1476 n1486 INVx1_ASAP7_75t_R
XU1859 n1478 n1487 INVx1_ASAP7_75t_R
XU1860 n1480 n1488 INVx1_ASAP7_75t_R
XU1861 n1489 add_6_root_r893_B_1_ INVx1_ASAP7_75t_R
XU1862 n1491 add_6_root_r893_B_2_ INVx1_ASAP7_75t_R
XU1863 n1493 add_6_root_r893_B_3_ INVx1_ASAP7_75t_R
XU1864 n1495 add_6_root_r893_B_4_ INVx1_ASAP7_75t_R
XU1865 n1497 add_6_root_r893_B_5_ INVx1_ASAP7_75t_R
XU1866 n1499 add_6_root_r893_B_6_ INVx1_ASAP7_75t_R
XU1867 n1501 add_6_root_r893_B_7_ INVx1_ASAP7_75t_R
XU1868 n1503 add_6_root_r893_B_8_ INVx1_ASAP7_75t_R
XU1869 n1504 add_6_root_r893_B_9_ INVx1_ASAP7_75t_R
XU1870 n1490 n1505 INVx1_ASAP7_75t_R
XU1871 n1492 n1506 INVx1_ASAP7_75t_R
XU1872 n1494 n1507 INVx1_ASAP7_75t_R
XU1873 n1496 n1508 INVx1_ASAP7_75t_R
XU1874 n1498 n1509 INVx1_ASAP7_75t_R
XU1875 n1500 n1510 INVx1_ASAP7_75t_R
XU1876 n1502 n1511 INVx1_ASAP7_75t_R
XU1877 n1512 N1246 INVx1_ASAP7_75t_R
XU1878 n1514 N1247 INVx1_ASAP7_75t_R
XU1879 n1516 N1248 INVx1_ASAP7_75t_R
XU1880 n1518 N1249 INVx1_ASAP7_75t_R
XU1881 n1520 N1250 INVx1_ASAP7_75t_R
XU1882 n1522 N1251 INVx1_ASAP7_75t_R
XU1883 n1524 N1252 INVx1_ASAP7_75t_R
XU1884 n1525 N1253 INVx1_ASAP7_75t_R
XU1885 n1513 n1526 INVx1_ASAP7_75t_R
XU1886 n1515 n1527 INVx1_ASAP7_75t_R
XU1887 n1517 n1528 INVx1_ASAP7_75t_R
XU1888 n1519 n1529 INVx1_ASAP7_75t_R
XU1889 n1521 n1530 INVx1_ASAP7_75t_R
XU1890 n1523 n1531 INVx1_ASAP7_75t_R
XU1891 n1532 N1099 INVx1_ASAP7_75t_R
XU1892 n1534 N1100 INVx1_ASAP7_75t_R
XU1893 n1536 N1101 INVx1_ASAP7_75t_R
XU1894 n1538 N1102 INVx1_ASAP7_75t_R
XU1895 n1540 N1103 INVx1_ASAP7_75t_R
XU1896 n1542 N1104 INVx1_ASAP7_75t_R
XU1897 n1544 N1105 INVx1_ASAP7_75t_R
XU1898 n1545 N1106 INVx1_ASAP7_75t_R
XU1899 n1533 n1546 INVx1_ASAP7_75t_R
XU1900 n1535 n1547 INVx1_ASAP7_75t_R
XU1901 n1537 n1548 INVx1_ASAP7_75t_R
XU1902 n1539 n1549 INVx1_ASAP7_75t_R
XU1903 n1541 n1550 INVx1_ASAP7_75t_R
XU1904 n1543 n1551 INVx1_ASAP7_75t_R
XU1905 n1552 N763 INVx1_ASAP7_75t_R
XU1906 n1554 N764 INVx1_ASAP7_75t_R
XU1907 n1556 N765 INVx1_ASAP7_75t_R
XU1908 n1558 N766 INVx1_ASAP7_75t_R
XU1909 n1560 N767 INVx1_ASAP7_75t_R
XU1910 n1562 N768 INVx1_ASAP7_75t_R
XU1911 n1564 N769 INVx1_ASAP7_75t_R
XU1912 n1566 N770 INVx1_ASAP7_75t_R
XU1913 n1567 N771 INVx1_ASAP7_75t_R
XU1914 n1553 n1568 INVx1_ASAP7_75t_R
XU1915 n1555 n1569 INVx1_ASAP7_75t_R
XU1916 n1557 n1570 INVx1_ASAP7_75t_R
XU1917 n1559 n1571 INVx1_ASAP7_75t_R
XU1918 n1561 n1572 INVx1_ASAP7_75t_R
XU1919 n1563 n1573 INVx1_ASAP7_75t_R
XU1920 n1565 n1574 INVx1_ASAP7_75t_R
XU1921 n1575 N1120 INVx1_ASAP7_75t_R
XU1922 n1577 N1121 INVx1_ASAP7_75t_R
XU1923 n1579 N1122 INVx1_ASAP7_75t_R
XU1924 n1581 N1123 INVx1_ASAP7_75t_R
XU1925 n1583 N1124 INVx1_ASAP7_75t_R
XU1926 n1585 N1125 INVx1_ASAP7_75t_R
XU1927 n1587 N1126 INVx1_ASAP7_75t_R
XU1928 n1588 N1127 INVx1_ASAP7_75t_R
XU1929 n1576 n1589 INVx1_ASAP7_75t_R
XU1930 n1578 n1590 INVx1_ASAP7_75t_R
XU1931 n1580 n1591 INVx1_ASAP7_75t_R
XU1932 n1582 n1592 INVx1_ASAP7_75t_R
XU1933 n1584 n1593 INVx1_ASAP7_75t_R
XU1934 n1586 n1594 INVx1_ASAP7_75t_R
XU1935 n1595 N1225 INVx1_ASAP7_75t_R
XU1936 n1597 N1226 INVx1_ASAP7_75t_R
XU1937 n1599 N1227 INVx1_ASAP7_75t_R
XU1938 n1601 N1228 INVx1_ASAP7_75t_R
XU1939 n1603 N1229 INVx1_ASAP7_75t_R
XU1940 n1605 N1230 INVx1_ASAP7_75t_R
XU1941 n1607 N1231 INVx1_ASAP7_75t_R
XU1942 n1608 N1232 INVx1_ASAP7_75t_R
XU1943 n1596 n1609 INVx1_ASAP7_75t_R
XU1944 n1598 n1610 INVx1_ASAP7_75t_R
XU1945 n1600 n1611 INVx1_ASAP7_75t_R
XU1946 n1602 n1612 INVx1_ASAP7_75t_R
XU1947 n1604 n1613 INVx1_ASAP7_75t_R
XU1948 n1606 n1614 INVx1_ASAP7_75t_R
XU1949 n1615 N784 INVx1_ASAP7_75t_R
XU1950 n1617 N785 INVx1_ASAP7_75t_R
XU1951 n1619 N786 INVx1_ASAP7_75t_R
XU1952 n1621 N787 INVx1_ASAP7_75t_R
XU1953 n1623 N788 INVx1_ASAP7_75t_R
XU1954 n1625 N789 INVx1_ASAP7_75t_R
XU1955 n1627 N790 INVx1_ASAP7_75t_R
XU1956 n1629 N791 INVx1_ASAP7_75t_R
XU1957 n1630 N792 INVx1_ASAP7_75t_R
XU1958 n1616 n1631 INVx1_ASAP7_75t_R
XU1959 n1618 n1632 INVx1_ASAP7_75t_R
XU1960 n1620 n1633 INVx1_ASAP7_75t_R
XU1961 n1622 n1634 INVx1_ASAP7_75t_R
XU1962 n1624 n1635 INVx1_ASAP7_75t_R
XU1963 n1626 n1636 INVx1_ASAP7_75t_R
XU1964 n1628 n1637 INVx1_ASAP7_75t_R
XU1965 n1638 N931 INVx1_ASAP7_75t_R
XU1966 n1640 N932 INVx1_ASAP7_75t_R
XU1967 n1642 N933 INVx1_ASAP7_75t_R
XU1968 n1644 N934 INVx1_ASAP7_75t_R
XU1969 n1646 N935 INVx1_ASAP7_75t_R
XU1970 n1648 N936 INVx1_ASAP7_75t_R
XU1971 n1650 N937 INVx1_ASAP7_75t_R
XU1972 n1651 N938 INVx1_ASAP7_75t_R
XU1973 n1639 n1652 INVx1_ASAP7_75t_R
XU1974 n1641 n1653 INVx1_ASAP7_75t_R
XU1975 n1643 n1654 INVx1_ASAP7_75t_R
XU1976 n1645 n1655 INVx1_ASAP7_75t_R
XU1977 n1647 n1656 INVx1_ASAP7_75t_R
XU1978 n1649 n1657 INVx1_ASAP7_75t_R
XU1979 n1658 N826 INVx1_ASAP7_75t_R
XU1980 n1660 N827 INVx1_ASAP7_75t_R
XU1981 n1662 N828 INVx1_ASAP7_75t_R
XU1982 n1664 N829 INVx1_ASAP7_75t_R
XU1983 n1666 N830 INVx1_ASAP7_75t_R
XU1984 n1668 N831 INVx1_ASAP7_75t_R
XU1985 n1670 N832 INVx1_ASAP7_75t_R
XU1986 n1671 N833 INVx1_ASAP7_75t_R
XU1987 n1659 n1672 INVx1_ASAP7_75t_R
XU1988 n1661 n1673 INVx1_ASAP7_75t_R
XU1989 n1663 n1674 INVx1_ASAP7_75t_R
XU1990 n1665 n1675 INVx1_ASAP7_75t_R
XU1991 n1667 n1676 INVx1_ASAP7_75t_R
XU1992 n1669 n1677 INVx1_ASAP7_75t_R
XU1993 n1678 N805 INVx1_ASAP7_75t_R
XU1994 n1680 N806 INVx1_ASAP7_75t_R
XU1995 n1682 N807 INVx1_ASAP7_75t_R
XU1996 n1684 N808 INVx1_ASAP7_75t_R
XU1997 n1686 N809 INVx1_ASAP7_75t_R
XU1998 n1688 N810 INVx1_ASAP7_75t_R
XU1999 n1690 N811 INVx1_ASAP7_75t_R
XU2000 n1692 N812 INVx1_ASAP7_75t_R
XU2001 n1693 N813 INVx1_ASAP7_75t_R
XU2002 n1679 n1694 INVx1_ASAP7_75t_R
XU2003 n1681 n1695 INVx1_ASAP7_75t_R
XU2004 n1683 n1696 INVx1_ASAP7_75t_R
XU2005 n1685 n1697 INVx1_ASAP7_75t_R
XU2006 n1687 n1698 INVx1_ASAP7_75t_R
XU2007 n1689 n1699 INVx1_ASAP7_75t_R
XU2008 n1691 n1700 INVx1_ASAP7_75t_R
XU2009 n1701 N847 INVx1_ASAP7_75t_R
XU2010 n1703 N848 INVx1_ASAP7_75t_R
XU2011 n1705 N849 INVx1_ASAP7_75t_R
XU2012 n1707 N850 INVx1_ASAP7_75t_R
XU2013 n1709 N851 INVx1_ASAP7_75t_R
XU2014 n1711 N852 INVx1_ASAP7_75t_R
XU2015 n1713 N853 INVx1_ASAP7_75t_R
XU2016 n1714 N854 INVx1_ASAP7_75t_R
XU2017 n1702 n1715 INVx1_ASAP7_75t_R
XU2018 n1704 n1716 INVx1_ASAP7_75t_R
XU2019 n1706 n1717 INVx1_ASAP7_75t_R
XU2020 n1708 n1718 INVx1_ASAP7_75t_R
XU2021 n1710 n1719 INVx1_ASAP7_75t_R
XU2022 n1712 n1720 INVx1_ASAP7_75t_R
XU2023 n1721 N868 INVx1_ASAP7_75t_R
XU2024 n1723 N869 INVx1_ASAP7_75t_R
XU2025 n1725 N870 INVx1_ASAP7_75t_R
XU2026 n1727 N871 INVx1_ASAP7_75t_R
XU2027 n1729 N872 INVx1_ASAP7_75t_R
XU2028 n1731 N873 INVx1_ASAP7_75t_R
XU2029 n1733 N874 INVx1_ASAP7_75t_R
XU2030 n1734 N875 INVx1_ASAP7_75t_R
XU2031 n1722 n1735 INVx1_ASAP7_75t_R
XU2032 n1724 n1736 INVx1_ASAP7_75t_R
XU2033 n1726 n1737 INVx1_ASAP7_75t_R
XU2034 n1728 n1738 INVx1_ASAP7_75t_R
XU2035 n1730 n1739 INVx1_ASAP7_75t_R
XU2036 n1732 n1740 INVx1_ASAP7_75t_R
XU2037 n1741 N889 INVx1_ASAP7_75t_R
XU2038 n1743 N890 INVx1_ASAP7_75t_R
XU2039 n1745 N891 INVx1_ASAP7_75t_R
XU2040 n1747 N892 INVx1_ASAP7_75t_R
XU2041 n1749 N893 INVx1_ASAP7_75t_R
XU2042 n1751 N894 INVx1_ASAP7_75t_R
XU2043 n1753 N895 INVx1_ASAP7_75t_R
XU2044 n1754 N896 INVx1_ASAP7_75t_R
XU2045 n1742 n1755 INVx1_ASAP7_75t_R
XU2046 n1744 n1756 INVx1_ASAP7_75t_R
XU2047 n1746 n1757 INVx1_ASAP7_75t_R
XU2048 n1748 n1758 INVx1_ASAP7_75t_R
XU2049 n1750 n1759 INVx1_ASAP7_75t_R
XU2050 n1752 n1760 INVx1_ASAP7_75t_R
XU2051 n1761 N973 INVx1_ASAP7_75t_R
XU2052 n1763 N974 INVx1_ASAP7_75t_R
XU2053 n1765 N975 INVx1_ASAP7_75t_R
XU2054 n1767 N976 INVx1_ASAP7_75t_R
XU2055 n1769 N977 INVx1_ASAP7_75t_R
XU2056 n1771 N978 INVx1_ASAP7_75t_R
XU2057 n1773 N979 INVx1_ASAP7_75t_R
XU2058 n1774 N980 INVx1_ASAP7_75t_R
XU2059 n1762 n1775 INVx1_ASAP7_75t_R
XU2060 n1764 n1776 INVx1_ASAP7_75t_R
XU2061 n1766 n1777 INVx1_ASAP7_75t_R
XU2062 n1768 n1778 INVx1_ASAP7_75t_R
XU2063 n1770 n1779 INVx1_ASAP7_75t_R
XU2064 n1772 n1780 INVx1_ASAP7_75t_R
XU2065 n1781 N1057 INVx1_ASAP7_75t_R
XU2066 n1783 N1058 INVx1_ASAP7_75t_R
XU2067 n1785 N1059 INVx1_ASAP7_75t_R
XU2068 n1787 N1060 INVx1_ASAP7_75t_R
XU2069 n1789 N1061 INVx1_ASAP7_75t_R
XU2070 n1791 N1062 INVx1_ASAP7_75t_R
XU2071 n1793 N1063 INVx1_ASAP7_75t_R
XU2072 n1795 N1064 INVx1_ASAP7_75t_R
XU2073 n1796 N1065 INVx1_ASAP7_75t_R
XU2074 n1782 n1797 INVx1_ASAP7_75t_R
XU2075 n1784 n1798 INVx1_ASAP7_75t_R
XU2076 n1786 n1799 INVx1_ASAP7_75t_R
XU2077 n1788 n1800 INVx1_ASAP7_75t_R
XU2078 n1790 n1801 INVx1_ASAP7_75t_R
XU2079 n1792 n1802 INVx1_ASAP7_75t_R
XU2080 n1794 n1803 INVx1_ASAP7_75t_R
XU2081 n1804 N1204 INVx1_ASAP7_75t_R
XU2082 n1806 N1205 INVx1_ASAP7_75t_R
XU2083 n1808 N1206 INVx1_ASAP7_75t_R
XU2084 n1810 N1207 INVx1_ASAP7_75t_R
XU2085 n1812 N1208 INVx1_ASAP7_75t_R
XU2086 n1814 N1209 INVx1_ASAP7_75t_R
XU2087 n1816 N1210 INVx1_ASAP7_75t_R
XU2088 n1818 N1211 INVx1_ASAP7_75t_R
XU2089 n1819 N1212 INVx1_ASAP7_75t_R
XU2090 n1805 n1820 INVx1_ASAP7_75t_R
XU2091 n1807 n1821 INVx1_ASAP7_75t_R
XU2092 n1809 n1822 INVx1_ASAP7_75t_R
XU2093 n1811 n1823 INVx1_ASAP7_75t_R
XU2094 n1813 n1824 INVx1_ASAP7_75t_R
XU2095 n1815 n1825 INVx1_ASAP7_75t_R
XU2096 n1817 n1826 INVx1_ASAP7_75t_R
XU2097 n1844 add_4_root_r893_SUM_10_ INVx1_ASAP7_75t_R
XU2098 n1827 add_4_root_r893_SUM_1_ INVx1_ASAP7_75t_R
XU2099 n1829 add_4_root_r893_SUM_2_ INVx1_ASAP7_75t_R
XU2100 n1831 add_4_root_r893_SUM_3_ INVx1_ASAP7_75t_R
XU2101 n1833 add_4_root_r893_SUM_4_ INVx1_ASAP7_75t_R
XU2102 n1835 add_4_root_r893_SUM_5_ INVx1_ASAP7_75t_R
XU2103 n1837 add_4_root_r893_SUM_6_ INVx1_ASAP7_75t_R
XU2104 n1839 add_4_root_r893_SUM_7_ INVx1_ASAP7_75t_R
XU2105 n1841 add_4_root_r893_SUM_8_ INVx1_ASAP7_75t_R
XU2106 n1843 add_4_root_r893_SUM_9_ INVx1_ASAP7_75t_R
XU2107 n1828 n1845 INVx1_ASAP7_75t_R
XU2108 n1830 n1846 INVx1_ASAP7_75t_R
XU2109 n1832 n1847 INVx1_ASAP7_75t_R
XU2110 n1834 n1848 INVx1_ASAP7_75t_R
XU2111 n1836 n1849 INVx1_ASAP7_75t_R
XU2112 n1838 n1850 INVx1_ASAP7_75t_R
XU2113 n1840 n1851 INVx1_ASAP7_75t_R
XU2114 n1842 n1852 INVx1_ASAP7_75t_R
XU2115 n1870 N1024 INVx1_ASAP7_75t_R
XU2116 n1853 N1015 INVx1_ASAP7_75t_R
XU2117 n1855 N1016 INVx1_ASAP7_75t_R
XU2118 n1857 N1017 INVx1_ASAP7_75t_R
XU2119 n1859 N1018 INVx1_ASAP7_75t_R
XU2120 n1861 N1019 INVx1_ASAP7_75t_R
XU2121 n1863 N1020 INVx1_ASAP7_75t_R
XU2122 n1865 N1021 INVx1_ASAP7_75t_R
XU2123 n1867 N1022 INVx1_ASAP7_75t_R
XU2124 n1869 N1023 INVx1_ASAP7_75t_R
XU2125 n1854 n1871 INVx1_ASAP7_75t_R
XU2126 n1856 n1872 INVx1_ASAP7_75t_R
XU2127 n1858 n1873 INVx1_ASAP7_75t_R
XU2128 n1860 n1874 INVx1_ASAP7_75t_R
XU2129 n1862 n1875 INVx1_ASAP7_75t_R
XU2130 n1864 n1876 INVx1_ASAP7_75t_R
XU2131 n1866 n1877 INVx1_ASAP7_75t_R
XU2132 n1868 n1878 INVx1_ASAP7_75t_R
XU2133 n1896 N1045 INVx1_ASAP7_75t_R
XU2134 n1879 N1036 INVx1_ASAP7_75t_R
XU2135 n1881 N1037 INVx1_ASAP7_75t_R
XU2136 n1883 N1038 INVx1_ASAP7_75t_R
XU2137 n1885 N1039 INVx1_ASAP7_75t_R
XU2138 n1887 N1040 INVx1_ASAP7_75t_R
XU2139 n1889 N1041 INVx1_ASAP7_75t_R
XU2140 n1891 N1042 INVx1_ASAP7_75t_R
XU2141 n1893 N1043 INVx1_ASAP7_75t_R
XU2142 n1895 N1044 INVx1_ASAP7_75t_R
XU2143 n1880 n1897 INVx1_ASAP7_75t_R
XU2144 n1882 n1898 INVx1_ASAP7_75t_R
XU2145 n1884 n1899 INVx1_ASAP7_75t_R
XU2146 n1886 n1900 INVx1_ASAP7_75t_R
XU2147 n1888 n1901 INVx1_ASAP7_75t_R
XU2148 n1890 n1902 INVx1_ASAP7_75t_R
XU2149 n1892 n1903 INVx1_ASAP7_75t_R
XU2150 n1894 n1904 INVx1_ASAP7_75t_R
XU2151 state_cs n1906 INVx1_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW01_add_0 A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[12] SUM[11] SUM[10] SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] CO
XU1_11 A[11] B[11] n3 n13 n14 FAx1_ASAP7_75t_R
XU1_10 A[10] B[10] n4 n15 n16 FAx1_ASAP7_75t_R
XU1_9 A[9] B[9] n5 n17 n18 FAx1_ASAP7_75t_R
XU1_8 A[8] B[8] n6 n19 n20 FAx1_ASAP7_75t_R
XU1_7 A[7] B[7] n7 n21 n22 FAx1_ASAP7_75t_R
XU1_6 A[6] B[6] n8 n23 n24 FAx1_ASAP7_75t_R
XU1_5 A[5] B[5] n9 n25 n26 FAx1_ASAP7_75t_R
XU1_4 A[4] B[4] n10 n27 n28 FAx1_ASAP7_75t_R
XU1_3 A[3] B[3] n11 n29 n30 FAx1_ASAP7_75t_R
XU1_2 A[2] B[2] n12 n31 n32 FAx1_ASAP7_75t_R
XU1_1 A[1] B[1] n1 n33 n34 FAx1_ASAP7_75t_R
XU1 A[0] B[0] n1 AND2x2_ASAP7_75t_R
XU2 B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU3 n15 n3 INVx1_ASAP7_75t_R
XU4 n17 n4 INVx1_ASAP7_75t_R
XU5 n19 n5 INVx1_ASAP7_75t_R
XU6 n21 n6 INVx1_ASAP7_75t_R
XU7 n23 n7 INVx1_ASAP7_75t_R
XU8 n25 n8 INVx1_ASAP7_75t_R
XU9 n27 n9 INVx1_ASAP7_75t_R
XU10 n29 n10 INVx1_ASAP7_75t_R
XU11 n31 n11 INVx1_ASAP7_75t_R
XU12 n33 n12 INVx1_ASAP7_75t_R
XU13 n18 SUM[9] INVx1_ASAP7_75t_R
XU14 n20 SUM[8] INVx1_ASAP7_75t_R
XU15 n22 SUM[7] INVx1_ASAP7_75t_R
XU16 n24 SUM[6] INVx1_ASAP7_75t_R
XU17 n26 SUM[5] INVx1_ASAP7_75t_R
XU18 n28 SUM[4] INVx1_ASAP7_75t_R
XU19 n30 SUM[3] INVx1_ASAP7_75t_R
XU20 n32 SUM[2] INVx1_ASAP7_75t_R
XU21 n34 SUM[1] INVx1_ASAP7_75t_R
XU22 n13 SUM[12] INVx1_ASAP7_75t_R
XU23 n14 SUM[11] INVx1_ASAP7_75t_R
XU24 n16 SUM[10] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW01_add_1 A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[12] SUM[11] SUM[10] SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] CO
XU1_10 A[10] B[10] n3 n12 n13 FAx1_ASAP7_75t_R
XU1_9 A[9] B[9] n4 n14 n15 FAx1_ASAP7_75t_R
XU1_8 A[8] B[8] n5 n16 n17 FAx1_ASAP7_75t_R
XU1_7 A[7] B[7] n6 n18 n19 FAx1_ASAP7_75t_R
XU1_6 A[6] B[6] n7 n20 n21 FAx1_ASAP7_75t_R
XU1_5 A[5] B[5] n8 n22 n23 FAx1_ASAP7_75t_R
XU1_4 A[4] B[4] n9 n24 n25 FAx1_ASAP7_75t_R
XU1_3 A[3] B[3] n10 n26 n27 FAx1_ASAP7_75t_R
XU1_2 A[2] B[2] n11 n28 n29 FAx1_ASAP7_75t_R
XU1_1 A[1] B[1] n2 n30 n31 FAx1_ASAP7_75t_R
XU1 B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU2 A[0] B[0] n2 AND2x2_ASAP7_75t_R
XU3 n14 n3 INVx1_ASAP7_75t_R
XU4 n16 n4 INVx1_ASAP7_75t_R
XU5 n18 n5 INVx1_ASAP7_75t_R
XU6 n20 n6 INVx1_ASAP7_75t_R
XU7 n22 n7 INVx1_ASAP7_75t_R
XU8 n24 n8 INVx1_ASAP7_75t_R
XU9 n26 n9 INVx1_ASAP7_75t_R
XU10 n28 n10 INVx1_ASAP7_75t_R
XU11 n30 n11 INVx1_ASAP7_75t_R
XU12 n15 SUM[9] INVx1_ASAP7_75t_R
XU13 n17 SUM[8] INVx1_ASAP7_75t_R
XU14 n19 SUM[7] INVx1_ASAP7_75t_R
XU15 n21 SUM[6] INVx1_ASAP7_75t_R
XU16 n23 SUM[5] INVx1_ASAP7_75t_R
XU17 n25 SUM[4] INVx1_ASAP7_75t_R
XU18 n27 SUM[3] INVx1_ASAP7_75t_R
XU19 n29 SUM[2] INVx1_ASAP7_75t_R
XU20 n31 SUM[1] INVx1_ASAP7_75t_R
XU21 n12 SUM[11] INVx1_ASAP7_75t_R
XU22 n13 SUM[10] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW01_add_2 A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[12] SUM[11] SUM[10] SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] CO
XU1_10 A[10] B[10] n3 n12 n13 FAx1_ASAP7_75t_R
XU1_9 A[9] B[9] n4 n14 n15 FAx1_ASAP7_75t_R
XU1_8 A[8] B[8] n5 n16 n17 FAx1_ASAP7_75t_R
XU1_7 A[7] B[7] n6 n18 n19 FAx1_ASAP7_75t_R
XU1_6 A[6] B[6] n7 n20 n21 FAx1_ASAP7_75t_R
XU1_5 A[5] B[5] n8 n22 n23 FAx1_ASAP7_75t_R
XU1_4 A[4] B[4] n9 n24 n25 FAx1_ASAP7_75t_R
XU1_3 A[3] B[3] n10 n26 n27 FAx1_ASAP7_75t_R
XU1_2 A[2] B[2] n11 n28 n29 FAx1_ASAP7_75t_R
XU1_1 A[1] B[1] n1 n30 n31 FAx1_ASAP7_75t_R
XU1 A[0] B[0] n1 AND2x2_ASAP7_75t_R
XU2 B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU3 n14 n3 INVx1_ASAP7_75t_R
XU4 n16 n4 INVx1_ASAP7_75t_R
XU5 n18 n5 INVx1_ASAP7_75t_R
XU6 n20 n6 INVx1_ASAP7_75t_R
XU7 n22 n7 INVx1_ASAP7_75t_R
XU8 n24 n8 INVx1_ASAP7_75t_R
XU9 n26 n9 INVx1_ASAP7_75t_R
XU10 n28 n10 INVx1_ASAP7_75t_R
XU11 n30 n11 INVx1_ASAP7_75t_R
XU12 n15 SUM[9] INVx1_ASAP7_75t_R
XU13 n17 SUM[8] INVx1_ASAP7_75t_R
XU14 n19 SUM[7] INVx1_ASAP7_75t_R
XU15 n21 SUM[6] INVx1_ASAP7_75t_R
XU16 n23 SUM[5] INVx1_ASAP7_75t_R
XU17 n25 SUM[4] INVx1_ASAP7_75t_R
XU18 n27 SUM[3] INVx1_ASAP7_75t_R
XU19 n29 SUM[2] INVx1_ASAP7_75t_R
XU20 n31 SUM[1] INVx1_ASAP7_75t_R
XU21 n12 SUM[11] INVx1_ASAP7_75t_R
XU22 n13 SUM[10] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_0 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_1 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_2 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_3 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_4 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_5 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_6 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_7 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_8 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_9 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_10 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_11 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_12 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_13 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_14 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_15 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_16 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_17 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_18 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_19 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_20 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_21 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_22 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_23 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_24 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_25 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_26 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_27 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_28 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_29 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_30 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT CIM_DW_mult_uns_31 a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 a[2] n83 INVx1_ASAP7_75t_R
XU71 n35 n84 INVx1_ASAP7_75t_R
XU72 a[0] n85 INVx1_ASAP7_75t_R
XU73 b[3] n86 INVx1_ASAP7_75t_R
XU74 b[0] n87 INVx1_ASAP7_75t_R
XU75 n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


